# Copyright (c) 1993 - 2019 ARM Limited. All Rights Reserved.
# Use of this Software is subject to the terms and conditions of the
# applicable license agreement with ARM Limited.

# PhyVGen V 8.3.0
# ARM Version r4p0
# Creation Date: Mon Nov 11 12:00:01 2019


# Memory Configuration:
# ~~~~~~~~~~~~~~~~~~~~~
#  -activity_factor 50 -atf off -back_biasing off -bits 19 -bmux on
# -bus_notation on -check_instname off -diodes on -drive 6 -ema on -frequency
# 1.0 -instname rf2_32x19_wm0 -left_bus_delim "[" -mux 2 -mvt BASE -name_case
# upper -pipeline off -power_gating off -power_type otc -pwr_gnd_rename
# vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -rcols 2 -redundancy off -retention on
# -right_bus_delim "]" -rrows 0 -ser none -site_def off -top_layer m5-m10
# -words 32 -wp_size 1 -write_mask off -write_thru off -corners
# ff_0p99v_0p99v_125c,ss_0p81v_0p81v_m40c,tt_0p90v_0p90v_25c
# 

VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO rf2_32x19_wm0
	FOREIGN rf2_32x19_wm0 0 0 ;
	SYMMETRY X Y ;
	SIZE 21.165 BY 100.94 ;
	CLASS BLOCK ;
	PIN AA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 32.87 0.25 32.97 ;
			LAYER	M2 ;
			RECT	0 32.87 0.25 32.97 ;
			LAYER	M3 ;
			RECT	0 32.87 0.25 32.97 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[0]

	PIN AA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 35.9 0.25 36 ;
			LAYER	M2 ;
			RECT	0 35.9 0.25 36 ;
			LAYER	M3 ;
			RECT	0 35.9 0.25 36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[1]

	PIN AA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 38.93 0.25 39.03 ;
			LAYER	M2 ;
			RECT	0 38.93 0.25 39.03 ;
			LAYER	M3 ;
			RECT	0 38.93 0.25 39.03 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[2]

	PIN AA[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 40.475 0.25 40.575 ;
			LAYER	M2 ;
			RECT	0 40.475 0.25 40.575 ;
			LAYER	M3 ;
			RECT	0 40.475 0.25 40.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[3]

	PIN AA[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.505 0.25 43.605 ;
			LAYER	M2 ;
			RECT	0 43.505 0.25 43.605 ;
			LAYER	M3 ;
			RECT	0 43.505 0.25 43.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[4]

	PIN AB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.785 0.25 65.885 ;
			LAYER	M2 ;
			RECT	0 65.785 0.25 65.885 ;
			LAYER	M3 ;
			RECT	0 65.785 0.25 65.885 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[0]

	PIN AB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.56 0.25 62.66 ;
			LAYER	M2 ;
			RECT	0 62.56 0.25 62.66 ;
			LAYER	M3 ;
			RECT	0 62.56 0.25 62.66 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[1]

	PIN AB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.725 0.25 59.825 ;
			LAYER	M2 ;
			RECT	0 59.725 0.25 59.825 ;
			LAYER	M3 ;
			RECT	0 59.725 0.25 59.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[2]

	PIN AB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 58.18 0.25 58.28 ;
			LAYER	M2 ;
			RECT	0 58.18 0.25 58.28 ;
			LAYER	M3 ;
			RECT	0 58.18 0.25 58.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[3]

	PIN AB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 55.15 0.25 55.25 ;
			LAYER	M2 ;
			RECT	0 55.15 0.25 55.25 ;
			LAYER	M3 ;
			RECT	0 55.15 0.25 55.25 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[4]

	PIN AYA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.275 0.25 33.375 ;
			LAYER	M2 ;
			RECT	0 33.275 0.25 33.375 ;
			LAYER	M3 ;
			RECT	0 33.275 0.25 33.375 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[0]

	PIN AYA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.305 0.25 36.405 ;
			LAYER	M2 ;
			RECT	0 36.305 0.25 36.405 ;
			LAYER	M3 ;
			RECT	0 36.305 0.25 36.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[1]

	PIN AYA[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.335 0.25 39.435 ;
			LAYER	M2 ;
			RECT	0 39.335 0.25 39.435 ;
			LAYER	M3 ;
			RECT	0 39.335 0.25 39.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[2]

	PIN AYA[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 40.1 0.25 40.2 ;
			LAYER	M2 ;
			RECT	0 40.1 0.25 40.2 ;
			LAYER	M3 ;
			RECT	0 40.1 0.25 40.2 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[3]

	PIN AYA[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.305 0.25 43.405 ;
			LAYER	M2 ;
			RECT	0 43.305 0.25 43.405 ;
			LAYER	M3 ;
			RECT	0 43.305 0.25 43.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[4]

	PIN AYB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.38 0.25 65.48 ;
			LAYER	M2 ;
			RECT	0 65.38 0.25 65.48 ;
			LAYER	M3 ;
			RECT	0 65.38 0.25 65.48 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[0]

	PIN AYB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.35 0.25 62.45 ;
			LAYER	M2 ;
			RECT	0 62.35 0.25 62.45 ;
			LAYER	M3 ;
			RECT	0 62.35 0.25 62.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[1]

	PIN AYB[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.35 0.25 59.45 ;
			LAYER	M2 ;
			RECT	0 59.35 0.25 59.45 ;
			LAYER	M3 ;
			RECT	0 59.35 0.25 59.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[2]

	PIN AYB[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 58.585 0.25 58.685 ;
			LAYER	M2 ;
			RECT	0 58.585 0.25 58.685 ;
			LAYER	M3 ;
			RECT	0 58.585 0.25 58.685 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[3]

	PIN AYB[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 55.525 0.25 55.625 ;
			LAYER	M2 ;
			RECT	0 55.525 0.25 55.625 ;
			LAYER	M3 ;
			RECT	0 55.525 0.25 55.625 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[4]

	PIN CENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.11 0.25 30.21 ;
			LAYER	M2 ;
			RECT	0 30.11 0.25 30.21 ;
			LAYER	M3 ;
			RECT	0 30.11 0.25 30.21 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENA

	PIN CENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 70.305 0.25 70.405 ;
			LAYER	M2 ;
			RECT	0 70.305 0.25 70.405 ;
			LAYER	M3 ;
			RECT	0 70.305 0.25 70.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENB

	PIN CENYA
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 28.7 0.25 28.8 ;
			LAYER	M2 ;
			RECT	0 28.7 0.25 28.8 ;
			LAYER	M3 ;
			RECT	0 28.7 0.25 28.8 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENYA

	PIN CENYB
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 70.85 0.25 70.95 ;
			LAYER	M2 ;
			RECT	0 70.85 0.25 70.95 ;
			LAYER	M3 ;
			RECT	0 70.85 0.25 70.95 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENYB

	PIN CLKA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.73 0.25 39.83 ;
			LAYER	M2 ;
			RECT	0 39.73 0.25 39.83 ;
			LAYER	M3 ;
			RECT	0 39.73 0.25 39.83 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CLKA

	PIN CLKB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.38 0.25 60.48 ;
			LAYER	M2 ;
			RECT	0 60.38 0.25 60.48 ;
			LAYER	M3 ;
			RECT	0 60.38 0.25 60.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CLKB

	PIN COLLDISN
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.9 0.25 48 ;
			LAYER	M2 ;
			RECT	0 47.9 0.25 48 ;
			LAYER	M3 ;
			RECT	0 47.9 0.25 48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END COLLDISN

	PIN DB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 2.195 0.25 2.295 ;
			LAYER	M2 ;
			RECT	0 2.195 0.25 2.295 ;
			LAYER	M3 ;
			RECT	0 2.195 0.25 2.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[0]

	PIN DB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 75.605 0.25 75.705 ;
			LAYER	M2 ;
			RECT	0 75.605 0.25 75.705 ;
			LAYER	M3 ;
			RECT	0 75.605 0.25 75.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[10]

	PIN DB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 78.485 0.25 78.585 ;
			LAYER	M2 ;
			RECT	0 78.485 0.25 78.585 ;
			LAYER	M3 ;
			RECT	0 78.485 0.25 78.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[11]

	PIN DB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 81.365 0.25 81.465 ;
			LAYER	M2 ;
			RECT	0 81.365 0.25 81.465 ;
			LAYER	M3 ;
			RECT	0 81.365 0.25 81.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[12]

	PIN DB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 84.245 0.25 84.345 ;
			LAYER	M2 ;
			RECT	0 84.245 0.25 84.345 ;
			LAYER	M3 ;
			RECT	0 84.245 0.25 84.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[13]

	PIN DB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 87.125 0.25 87.225 ;
			LAYER	M2 ;
			RECT	0 87.125 0.25 87.225 ;
			LAYER	M3 ;
			RECT	0 87.125 0.25 87.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[14]

	PIN DB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 90.005 0.25 90.105 ;
			LAYER	M2 ;
			RECT	0 90.005 0.25 90.105 ;
			LAYER	M3 ;
			RECT	0 90.005 0.25 90.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[15]

	PIN DB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 92.885 0.25 92.985 ;
			LAYER	M2 ;
			RECT	0 92.885 0.25 92.985 ;
			LAYER	M3 ;
			RECT	0 92.885 0.25 92.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[16]

	PIN DB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 95.765 0.25 95.865 ;
			LAYER	M2 ;
			RECT	0 95.765 0.25 95.865 ;
			LAYER	M3 ;
			RECT	0 95.765 0.25 95.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[17]

	PIN DB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 98.645 0.25 98.745 ;
			LAYER	M2 ;
			RECT	0 98.645 0.25 98.745 ;
			LAYER	M3 ;
			RECT	0 98.645 0.25 98.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[18]

	PIN DB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 5.075 0.25 5.175 ;
			LAYER	M2 ;
			RECT	0 5.075 0.25 5.175 ;
			LAYER	M3 ;
			RECT	0 5.075 0.25 5.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[1]

	PIN DB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.955 0.25 8.055 ;
			LAYER	M2 ;
			RECT	0 7.955 0.25 8.055 ;
			LAYER	M3 ;
			RECT	0 7.955 0.25 8.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[2]

	PIN DB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.835 0.25 10.935 ;
			LAYER	M2 ;
			RECT	0 10.835 0.25 10.935 ;
			LAYER	M3 ;
			RECT	0 10.835 0.25 10.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[3]

	PIN DB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.715 0.25 13.815 ;
			LAYER	M2 ;
			RECT	0 13.715 0.25 13.815 ;
			LAYER	M3 ;
			RECT	0 13.715 0.25 13.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[4]

	PIN DB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.595 0.25 16.695 ;
			LAYER	M2 ;
			RECT	0 16.595 0.25 16.695 ;
			LAYER	M3 ;
			RECT	0 16.595 0.25 16.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[5]

	PIN DB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.475 0.25 19.575 ;
			LAYER	M2 ;
			RECT	0 19.475 0.25 19.575 ;
			LAYER	M3 ;
			RECT	0 19.475 0.25 19.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[6]

	PIN DB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.355 0.25 22.455 ;
			LAYER	M2 ;
			RECT	0 22.355 0.25 22.455 ;
			LAYER	M3 ;
			RECT	0 22.355 0.25 22.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[7]

	PIN DB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.235 0.25 25.335 ;
			LAYER	M2 ;
			RECT	0 25.235 0.25 25.335 ;
			LAYER	M3 ;
			RECT	0 25.235 0.25 25.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[8]

	PIN DB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 72.725 0.25 72.825 ;
			LAYER	M2 ;
			RECT	0 72.725 0.25 72.825 ;
			LAYER	M3 ;
			RECT	0 72.725 0.25 72.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[9]

	PIN DFTRAMBYP
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 67.3 0.25 67.4 ;
			LAYER	M2 ;
			RECT	0 67.3 0.25 67.4 ;
			LAYER	M3 ;
			RECT	0 67.3 0.25 67.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DFTRAMBYP

	PIN EMAA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 41.37 0.25 41.47 ;
			LAYER	M2 ;
			RECT	0 41.37 0.25 41.47 ;
			LAYER	M3 ;
			RECT	0 41.37 0.25 41.47 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[0]

	PIN EMAA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 41.17 0.25 41.27 ;
			LAYER	M2 ;
			RECT	0 41.17 0.25 41.27 ;
			LAYER	M3 ;
			RECT	0 41.17 0.25 41.27 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[1]

	PIN EMAA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.105 0.25 43.205 ;
			LAYER	M2 ;
			RECT	0 43.105 0.25 43.205 ;
			LAYER	M3 ;
			RECT	0 43.105 0.25 43.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[2]

	PIN EMAB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 55.905 0.25 56.005 ;
			LAYER	M2 ;
			RECT	0 55.905 0.25 56.005 ;
			LAYER	M3 ;
			RECT	0 55.905 0.25 56.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[0]

	PIN EMAB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.905 0.25 57.005 ;
			LAYER	M2 ;
			RECT	0 56.905 0.25 57.005 ;
			LAYER	M3 ;
			RECT	0 56.905 0.25 57.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[1]

	PIN EMAB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.425 0.25 54.525 ;
			LAYER	M2 ;
			RECT	0 54.425 0.25 54.525 ;
			LAYER	M3 ;
			RECT	0 54.425 0.25 54.525 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[2]

	PIN EMASA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 29.05 0.25 29.15 ;
			LAYER	M2 ;
			RECT	0 29.05 0.25 29.15 ;
			LAYER	M3 ;
			RECT	0 29.05 0.25 29.15 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMASA

	PIN QA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 2.455 0.25 2.555 ;
			LAYER	M2 ;
			RECT	0 2.455 0.25 2.555 ;
			LAYER	M3 ;
			RECT	0 2.455 0.25 2.555 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[0]

	PIN QA[10]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 75.345 0.25 75.445 ;
			LAYER	M2 ;
			RECT	0 75.345 0.25 75.445 ;
			LAYER	M3 ;
			RECT	0 75.345 0.25 75.445 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[10]

	PIN QA[11]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 78.225 0.25 78.325 ;
			LAYER	M2 ;
			RECT	0 78.225 0.25 78.325 ;
			LAYER	M3 ;
			RECT	0 78.225 0.25 78.325 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[11]

	PIN QA[12]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 81.105 0.25 81.205 ;
			LAYER	M2 ;
			RECT	0 81.105 0.25 81.205 ;
			LAYER	M3 ;
			RECT	0 81.105 0.25 81.205 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[12]

	PIN QA[13]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 83.985 0.25 84.085 ;
			LAYER	M2 ;
			RECT	0 83.985 0.25 84.085 ;
			LAYER	M3 ;
			RECT	0 83.985 0.25 84.085 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[13]

	PIN QA[14]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 86.865 0.25 86.965 ;
			LAYER	M2 ;
			RECT	0 86.865 0.25 86.965 ;
			LAYER	M3 ;
			RECT	0 86.865 0.25 86.965 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[14]

	PIN QA[15]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 89.745 0.25 89.845 ;
			LAYER	M2 ;
			RECT	0 89.745 0.25 89.845 ;
			LAYER	M3 ;
			RECT	0 89.745 0.25 89.845 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[15]

	PIN QA[16]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 92.625 0.25 92.725 ;
			LAYER	M2 ;
			RECT	0 92.625 0.25 92.725 ;
			LAYER	M3 ;
			RECT	0 92.625 0.25 92.725 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[16]

	PIN QA[17]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 95.505 0.25 95.605 ;
			LAYER	M2 ;
			RECT	0 95.505 0.25 95.605 ;
			LAYER	M3 ;
			RECT	0 95.505 0.25 95.605 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[17]

	PIN QA[18]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 98.385 0.25 98.485 ;
			LAYER	M2 ;
			RECT	0 98.385 0.25 98.485 ;
			LAYER	M3 ;
			RECT	0 98.385 0.25 98.485 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[18]

	PIN QA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 5.335 0.25 5.435 ;
			LAYER	M2 ;
			RECT	0 5.335 0.25 5.435 ;
			LAYER	M3 ;
			RECT	0 5.335 0.25 5.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[1]

	PIN QA[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 8.215 0.25 8.315 ;
			LAYER	M2 ;
			RECT	0 8.215 0.25 8.315 ;
			LAYER	M3 ;
			RECT	0 8.215 0.25 8.315 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[2]

	PIN QA[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 11.095 0.25 11.195 ;
			LAYER	M2 ;
			RECT	0 11.095 0.25 11.195 ;
			LAYER	M3 ;
			RECT	0 11.095 0.25 11.195 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[3]

	PIN QA[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.975 0.25 14.075 ;
			LAYER	M2 ;
			RECT	0 13.975 0.25 14.075 ;
			LAYER	M3 ;
			RECT	0 13.975 0.25 14.075 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[4]

	PIN QA[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.855 0.25 16.955 ;
			LAYER	M2 ;
			RECT	0 16.855 0.25 16.955 ;
			LAYER	M3 ;
			RECT	0 16.855 0.25 16.955 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[5]

	PIN QA[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.735 0.25 19.835 ;
			LAYER	M2 ;
			RECT	0 19.735 0.25 19.835 ;
			LAYER	M3 ;
			RECT	0 19.735 0.25 19.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[6]

	PIN QA[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.615 0.25 22.715 ;
			LAYER	M2 ;
			RECT	0 22.615 0.25 22.715 ;
			LAYER	M3 ;
			RECT	0 22.615 0.25 22.715 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[7]

	PIN QA[8]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.495 0.25 25.595 ;
			LAYER	M2 ;
			RECT	0 25.495 0.25 25.595 ;
			LAYER	M3 ;
			RECT	0 25.495 0.25 25.595 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[8]

	PIN QA[9]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 72.465 0.25 72.565 ;
			LAYER	M2 ;
			RECT	0 72.465 0.25 72.565 ;
			LAYER	M3 ;
			RECT	0 72.465 0.25 72.565 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[9]

	PIN RET1N
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 29.71 0.25 29.81 ;
			LAYER	M2 ;
			RECT	0 29.71 0.25 29.81 ;
			LAYER	M3 ;
			RECT	0 29.71 0.25 29.81 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END RET1N

	PIN SEA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.5 0.25 47.6 ;
			LAYER	M2 ;
			RECT	0 47.5 0.25 47.6 ;
			LAYER	M3 ;
			RECT	0 47.5 0.25 47.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SEA

	PIN SEB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 50.335 0.25 50.435 ;
			LAYER	M2 ;
			RECT	0 50.335 0.25 50.435 ;
			LAYER	M3 ;
			RECT	0 50.335 0.25 50.435 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SEB

	PIN SIA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.7 0.25 47.8 ;
			LAYER	M2 ;
			RECT	0 47.7 0.25 47.8 ;
			LAYER	M3 ;
			RECT	0 47.7 0.25 47.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIA[0]

	PIN SIA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 48.67 0.25 48.77 ;
			LAYER	M2 ;
			RECT	0 48.67 0.25 48.77 ;
			LAYER	M3 ;
			RECT	0 48.67 0.25 48.77 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIA[1]

	PIN SIB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 44.275 0.25 44.375 ;
			LAYER	M2 ;
			RECT	0 44.275 0.25 44.375 ;
			LAYER	M3 ;
			RECT	0 44.275 0.25 44.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIB[0]

	PIN SIB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 61.925 0.25 62.025 ;
			LAYER	M2 ;
			RECT	0 61.925 0.25 62.025 ;
			LAYER	M3 ;
			RECT	0 61.925 0.25 62.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIB[1]

	PIN SOA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 0.36 0.25 0.46 ;
			LAYER	M2 ;
			RECT	0 0.36 0.25 0.46 ;
			LAYER	M3 ;
			RECT	0 0.36 0.25 0.46 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOA[0]

	PIN SOA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 100.48 0.25 100.58 ;
			LAYER	M2 ;
			RECT	0 100.48 0.25 100.58 ;
			LAYER	M3 ;
			RECT	0 100.48 0.25 100.58 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOA[1]

	PIN SOB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 0.09 0.25 0.19 ;
			LAYER	M2 ;
			RECT	0 0.09 0.25 0.19 ;
			LAYER	M3 ;
			RECT	0 0.09 0.25 0.19 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOB[0]

	PIN SOB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 100.75 0.25 100.85 ;
			LAYER	M2 ;
			RECT	0 100.75 0.25 100.85 ;
			LAYER	M3 ;
			RECT	0 100.75 0.25 100.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOB[1]

	PIN TAA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 32.355 0.25 32.455 ;
			LAYER	M2 ;
			RECT	0 32.355 0.25 32.455 ;
			LAYER	M3 ;
			RECT	0 32.355 0.25 32.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[0]

	PIN TAA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 35.385 0.25 35.485 ;
			LAYER	M2 ;
			RECT	0 35.385 0.25 35.485 ;
			LAYER	M3 ;
			RECT	0 35.385 0.25 35.485 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[1]

	PIN TAA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 38.445 0.25 38.545 ;
			LAYER	M2 ;
			RECT	0 38.445 0.25 38.545 ;
			LAYER	M3 ;
			RECT	0 38.445 0.25 38.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[2]

	PIN TAA[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 40.96 0.25 41.06 ;
			LAYER	M2 ;
			RECT	0 40.96 0.25 41.06 ;
			LAYER	M3 ;
			RECT	0 40.96 0.25 41.06 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[3]

	PIN TAA[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.99 0.25 44.09 ;
			LAYER	M2 ;
			RECT	0 43.99 0.25 44.09 ;
			LAYER	M3 ;
			RECT	0 43.99 0.25 44.09 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[4]

	PIN TAB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 66.27 0.25 66.37 ;
			LAYER	M2 ;
			RECT	0 66.27 0.25 66.37 ;
			LAYER	M3 ;
			RECT	0 66.27 0.25 66.37 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[0]

	PIN TAB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 63.24 0.25 63.34 ;
			LAYER	M2 ;
			RECT	0 63.24 0.25 63.34 ;
			LAYER	M3 ;
			RECT	0 63.24 0.25 63.34 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[1]

	PIN TAB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.18 0.25 60.28 ;
			LAYER	M2 ;
			RECT	0 60.18 0.25 60.28 ;
			LAYER	M3 ;
			RECT	0 60.18 0.25 60.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[2]

	PIN TAB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 57.695 0.25 57.795 ;
			LAYER	M2 ;
			RECT	0 57.695 0.25 57.795 ;
			LAYER	M3 ;
			RECT	0 57.695 0.25 57.795 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[3]

	PIN TAB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.66 0.25 54.76 ;
			LAYER	M2 ;
			RECT	0 54.66 0.25 54.76 ;
			LAYER	M3 ;
			RECT	0 54.66 0.25 54.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[4]

	PIN TCENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 29.91 0.25 30.01 ;
			LAYER	M2 ;
			RECT	0 29.91 0.25 30.01 ;
			LAYER	M3 ;
			RECT	0 29.91 0.25 30.01 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TCENA

	PIN TCENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 69.91 0.25 70.01 ;
			LAYER	M2 ;
			RECT	0 69.91 0.25 70.01 ;
			LAYER	M3 ;
			RECT	0 69.91 0.25 70.01 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TCENB

	PIN TDB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 1.465 0.25 1.565 ;
			LAYER	M2 ;
			RECT	0 1.465 0.25 1.565 ;
			LAYER	M3 ;
			RECT	0 1.465 0.25 1.565 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[0]

	PIN TDB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 76.335 0.25 76.435 ;
			LAYER	M2 ;
			RECT	0 76.335 0.25 76.435 ;
			LAYER	M3 ;
			RECT	0 76.335 0.25 76.435 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[10]

	PIN TDB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.215 0.25 79.315 ;
			LAYER	M2 ;
			RECT	0 79.215 0.25 79.315 ;
			LAYER	M3 ;
			RECT	0 79.215 0.25 79.315 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[11]

	PIN TDB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.095 0.25 82.195 ;
			LAYER	M2 ;
			RECT	0 82.095 0.25 82.195 ;
			LAYER	M3 ;
			RECT	0 82.095 0.25 82.195 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[12]

	PIN TDB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 84.975 0.25 85.075 ;
			LAYER	M2 ;
			RECT	0 84.975 0.25 85.075 ;
			LAYER	M3 ;
			RECT	0 84.975 0.25 85.075 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[13]

	PIN TDB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 87.855 0.25 87.955 ;
			LAYER	M2 ;
			RECT	0 87.855 0.25 87.955 ;
			LAYER	M3 ;
			RECT	0 87.855 0.25 87.955 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[14]

	PIN TDB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 90.735 0.25 90.835 ;
			LAYER	M2 ;
			RECT	0 90.735 0.25 90.835 ;
			LAYER	M3 ;
			RECT	0 90.735 0.25 90.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[15]

	PIN TDB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 93.615 0.25 93.715 ;
			LAYER	M2 ;
			RECT	0 93.615 0.25 93.715 ;
			LAYER	M3 ;
			RECT	0 93.615 0.25 93.715 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[16]

	PIN TDB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 96.495 0.25 96.595 ;
			LAYER	M2 ;
			RECT	0 96.495 0.25 96.595 ;
			LAYER	M3 ;
			RECT	0 96.495 0.25 96.595 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[17]

	PIN TDB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 99.375 0.25 99.475 ;
			LAYER	M2 ;
			RECT	0 99.375 0.25 99.475 ;
			LAYER	M3 ;
			RECT	0 99.375 0.25 99.475 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[18]

	PIN TDB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 4.345 0.25 4.445 ;
			LAYER	M2 ;
			RECT	0 4.345 0.25 4.445 ;
			LAYER	M3 ;
			RECT	0 4.345 0.25 4.445 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[1]

	PIN TDB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.225 0.25 7.325 ;
			LAYER	M2 ;
			RECT	0 7.225 0.25 7.325 ;
			LAYER	M3 ;
			RECT	0 7.225 0.25 7.325 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[2]

	PIN TDB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.105 0.25 10.205 ;
			LAYER	M2 ;
			RECT	0 10.105 0.25 10.205 ;
			LAYER	M3 ;
			RECT	0 10.105 0.25 10.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[3]

	PIN TDB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 12.985 0.25 13.085 ;
			LAYER	M2 ;
			RECT	0 12.985 0.25 13.085 ;
			LAYER	M3 ;
			RECT	0 12.985 0.25 13.085 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[4]

	PIN TDB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 15.865 0.25 15.965 ;
			LAYER	M2 ;
			RECT	0 15.865 0.25 15.965 ;
			LAYER	M3 ;
			RECT	0 15.865 0.25 15.965 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[5]

	PIN TDB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 18.745 0.25 18.845 ;
			LAYER	M2 ;
			RECT	0 18.745 0.25 18.845 ;
			LAYER	M3 ;
			RECT	0 18.745 0.25 18.845 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[6]

	PIN TDB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 21.625 0.25 21.725 ;
			LAYER	M2 ;
			RECT	0 21.625 0.25 21.725 ;
			LAYER	M3 ;
			RECT	0 21.625 0.25 21.725 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[7]

	PIN TDB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 24.505 0.25 24.605 ;
			LAYER	M2 ;
			RECT	0 24.505 0.25 24.605 ;
			LAYER	M3 ;
			RECT	0 24.505 0.25 24.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[8]

	PIN TDB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 73.455 0.25 73.555 ;
			LAYER	M2 ;
			RECT	0 73.455 0.25 73.555 ;
			LAYER	M3 ;
			RECT	0 73.455 0.25 73.555 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[9]

	PIN TENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 32.05 0.25 32.15 ;
			LAYER	M2 ;
			RECT	0 32.05 0.25 32.15 ;
			LAYER	M3 ;
			RECT	0 32.05 0.25 32.15 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TENA

	PIN TENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 66.525 0.25 66.625 ;
			LAYER	M2 ;
			RECT	0 66.525 0.25 66.625 ;
			LAYER	M3 ;
			RECT	0 66.525 0.25 66.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TENB

	PIN VDDCE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 97.495 21.165 97.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 94.615 21.165 94.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 91.735 21.165 91.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 88.855 21.165 89.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 85.975 21.165 86.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 83.095 21.165 83.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 80.215 21.165 80.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 77.335 21.165 77.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 74.455 21.165 74.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 71.575 21.165 71.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.335 21.165 26.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.455 21.165 23.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 20.575 21.165 20.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 17.695 21.165 17.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 14.815 21.165 14.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 11.935 21.165 12.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.055 21.165 9.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.175 21.165 6.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.295 21.165 3.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.98 21.165 33.17 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 33.96 21.165 34.15 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 36.915 21.165 37.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 40.85 21.165 41.04 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 41.835 21.165 42.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 44.785 21.165 44.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 48.72 21.165 48.91 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.215 21.165 49.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 53.15 21.165 53.34 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 56.105 21.165 56.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 57.085 21.165 57.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.025 21.165 61.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 63.975 21.165 64.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.925 21.165 65.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 100.375 21.165 100.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.415 21.165 0.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 28.695 21.165 28.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.215 21.165 69.365 ;
		END

	END VDDCE

	PIN VDDPE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 99.915 21.165 100.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 97.035 21.165 97.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 94.155 21.165 94.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 91.275 21.165 91.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 88.395 21.165 88.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 85.515 21.165 85.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 82.635 21.165 82.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 79.755 21.165 79.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 76.875 21.165 77.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 73.995 21.165 74.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.915 21.165 24.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 21.035 21.165 21.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 18.155 21.165 18.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.275 21.165 15.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.395 21.165 12.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.515 21.165 9.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.635 21.165 6.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.755 21.165 3.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.875 21.165 1.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 30.025 21.165 30.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.03 21.165 32.22 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 34.945 21.165 35.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 35.93 21.165 36.12 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 37.9 21.165 38.09 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.88 21.165 39.07 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 39.865 21.165 40.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 42.82 21.165 43.01 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 46.755 21.165 46.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 47.74 21.165 47.93 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 50.2 21.165 50.39 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 51.18 21.165 51.37 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.12 21.165 55.31 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.07 21.165 58.26 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 59.055 21.165 59.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 60.04 21.165 60.23 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 62.005 21.165 62.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 62.99 21.165 63.18 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 65.91 21.165 66.1 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 67.91 21.165 68.1 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 100.605 21.165 100.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.185 21.165 0.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 28.235 21.165 28.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.675 21.165 69.825 ;
		END

	END VDDPE

	PIN VSSE
		USE GROUND ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 100.145 21.165 100.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.645 21.165 0.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 28.465 21.165 28.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.445 21.165 69.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 97.265 21.165 97.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 94.385 21.165 94.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.565 21.165 26.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.685 21.165 23.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 20.805 21.165 20.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 17.925 21.165 18.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.045 21.165 15.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.165 21.165 12.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.285 21.165 9.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.405 21.165 6.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 91.505 21.165 91.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.525 21.165 3.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 88.625 21.165 88.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 85.745 21.165 85.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 82.865 21.165 83.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 79.985 21.165 80.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 77.105 21.165 77.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 74.225 21.165 74.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 71.345 21.165 71.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 99.685 21.165 99.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 24.145 21.165 24.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 21.265 21.165 21.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 18.385 21.165 18.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 93.925 21.165 94.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.505 21.165 15.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.625 21.165 12.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.745 21.165 9.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.865 21.165 7.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.985 21.165 4.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 1.105 21.165 1.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 91.045 21.165 91.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 88.165 21.165 88.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 85.285 21.165 85.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 82.405 21.165 82.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 79.525 21.165 79.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 76.645 21.165 76.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 73.765 21.165 73.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 96.805 21.165 96.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.535 21.165 29.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 30.515 21.165 30.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.485 21.165 32.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 33.47 21.165 33.66 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 36.425 21.165 36.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 37.405 21.165 37.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.39 21.165 38.58 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 40.36 21.165 40.55 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 41.33 21.165 41.54 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 42.325 21.165 42.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 44.3 21.165 44.49 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 45.28 21.165 45.47 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 48.23 21.165 48.42 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.705 21.165 49.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.655 21.165 52.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 53.645 21.165 53.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.61 21.165 55.8 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 56.585 21.165 56.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 57.58 21.165 57.77 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 59.545 21.165 59.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 60.53 21.165 60.72 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.515 21.165 61.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.455 21.165 64.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 65.45 21.165 65.64 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 67.42 21.165 67.61 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 68.405 21.165 68.595 ;
		END

	END VSSE

	OBS
		LAYER	M1 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 20.845 100.59 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 1.665 0.32 2.095 ;
		RECT	0 2.655 0.32 4.245 ;
		RECT	0 4.545 0.32 4.975 ;
		RECT	0 5.535 0.32 7.125 ;
		RECT	0 7.425 0.32 7.855 ;
		RECT	0 8.415 0.32 10.005 ;
		RECT	0 10.305 0.32 10.735 ;
		RECT	0 11.295 0.32 12.885 ;
		RECT	0 13.185 0.32 13.615 ;
		RECT	0 14.175 0.32 15.765 ;
		RECT	0 16.065 0.32 16.495 ;
		RECT	0 17.055 0.32 18.645 ;
		RECT	0 18.945 0.32 19.375 ;
		RECT	0 19.935 0.32 21.525 ;
		RECT	0 21.825 0.32 22.255 ;
		RECT	0 22.815 0.32 24.405 ;
		RECT	0 24.705 0.32 25.135 ;
		RECT	0 25.695 0.32 28.6 ;
		RECT	0 28.9 0.32 28.95 ;
		RECT	0 29.25 0.32 29.61 ;
		RECT	0 30.31 0.32 31.95 ;
		RECT	0 32.555 0.32 32.77 ;
		RECT	0 33.07 0.32 33.175 ;
		RECT	0 33.475 0.32 35.285 ;
		RECT	0 35.585 0.32 35.8 ;
		RECT	0 36.1 0.32 36.205 ;
		RECT	0 36.505 0.32 38.345 ;
		RECT	0 38.645 0.32 38.83 ;
		RECT	0 39.13 0.32 39.235 ;
		RECT	0 39.535 0.32 39.63 ;
		RECT	0 39.93 0.32 40 ;
		RECT	0 40.3 0.32 40.375 ;
		RECT	0 40.675 0.32 40.86 ;
		RECT	0 41.57 0.32 43.005 ;
		RECT	0 43.705 0.32 43.89 ;
		RECT	0 44.475 0.32 47.4 ;
		RECT	0 48.1 0.32 48.57 ;
		RECT	0 48.87 0.32 50.235 ;
		RECT	0 50.535 0.32 54.325 ;
		RECT	0 54.86 0.32 55.05 ;
		RECT	0 55.35 0.32 55.425 ;
		RECT	0 55.725 0.32 55.805 ;
		RECT	0 56.105 0.32 56.805 ;
		RECT	0 57.105 0.32 57.595 ;
		RECT	0 57.895 0.32 58.08 ;
		RECT	0 58.38 0.32 58.485 ;
		RECT	0 58.785 0.32 59.25 ;
		RECT	0 59.55 0.32 59.625 ;
		RECT	0 59.925 0.32 60.08 ;
		RECT	0 60.58 0.32 61.825 ;
		RECT	0 62.125 0.32 62.25 ;
		RECT	0 62.76 0.32 63.14 ;
		RECT	0 63.44 0.32 65.28 ;
		RECT	0 65.58 0.32 65.685 ;
		RECT	0 65.985 0.32 66.17 ;
		RECT	0 66.725 0.32 67.2 ;
		RECT	0 67.5 0.32 69.81 ;
		RECT	0 70.11 0.32 70.205 ;
		RECT	0 70.505 0.32 70.75 ;
		RECT	0 71.05 0.32 72.365 ;
		RECT	0 72.925 0.32 73.355 ;
		RECT	0 73.655 0.32 75.245 ;
		RECT	0 75.805 0.32 76.235 ;
		RECT	0 76.535 0.32 78.125 ;
		RECT	0 78.685 0.32 79.115 ;
		RECT	0 79.415 0.32 81.005 ;
		RECT	0 81.565 0.32 81.995 ;
		RECT	0 82.295 0.32 83.885 ;
		RECT	0 84.445 0.32 84.875 ;
		RECT	0 85.175 0.32 86.765 ;
		RECT	0 87.325 0.32 87.755 ;
		RECT	0 88.055 0.32 89.645 ;
		RECT	0 90.205 0.32 90.635 ;
		RECT	0 90.935 0.32 92.525 ;
		RECT	0 93.085 0.32 93.515 ;
		RECT	0 93.815 0.32 95.405 ;
		RECT	0 95.965 0.32 96.395 ;
		RECT	0 96.695 0.32 98.285 ;
		RECT	0 98.845 0.32 99.275 ;
		RECT	0 99.575 0.32 100.38 ;
		RECT	20.845 0 21.165 100.94 ;
		RECT	0.32 0 20.845 0.35 ;
		RECT	0.32 100.59 20.845 100.94 ;
		LAYER	M2 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 20.845 100.59 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 1.665 0.32 2.095 ;
		RECT	0 2.655 0.32 4.245 ;
		RECT	0 4.545 0.32 4.975 ;
		RECT	0 5.535 0.32 7.125 ;
		RECT	0 7.425 0.32 7.855 ;
		RECT	0 8.415 0.32 10.005 ;
		RECT	0 10.305 0.32 10.735 ;
		RECT	0 11.295 0.32 12.885 ;
		RECT	0 13.185 0.32 13.615 ;
		RECT	0 14.175 0.32 15.765 ;
		RECT	0 16.065 0.32 16.495 ;
		RECT	0 17.055 0.32 18.645 ;
		RECT	0 18.945 0.32 19.375 ;
		RECT	0 19.935 0.32 21.525 ;
		RECT	0 21.825 0.32 22.255 ;
		RECT	0 22.815 0.32 24.405 ;
		RECT	0 24.705 0.32 25.135 ;
		RECT	0 25.695 0.32 28.6 ;
		RECT	0 28.9 0.32 28.95 ;
		RECT	0 29.25 0.32 29.61 ;
		RECT	0 30.31 0.32 31.95 ;
		RECT	0 32.555 0.32 32.77 ;
		RECT	0 33.07 0.32 33.175 ;
		RECT	0 33.475 0.32 35.285 ;
		RECT	0 35.585 0.32 35.8 ;
		RECT	0 36.1 0.32 36.205 ;
		RECT	0 36.505 0.32 38.345 ;
		RECT	0 38.645 0.32 38.83 ;
		RECT	0 39.13 0.32 39.235 ;
		RECT	0 39.535 0.32 39.63 ;
		RECT	0 39.93 0.32 40 ;
		RECT	0 40.3 0.32 40.375 ;
		RECT	0 40.675 0.32 40.86 ;
		RECT	0 41.57 0.32 43.005 ;
		RECT	0 43.705 0.32 43.89 ;
		RECT	0 44.475 0.32 47.4 ;
		RECT	0 48.1 0.32 48.57 ;
		RECT	0 48.87 0.32 50.235 ;
		RECT	0 50.535 0.32 54.325 ;
		RECT	0 54.86 0.32 55.05 ;
		RECT	0 55.35 0.32 55.425 ;
		RECT	0 55.725 0.32 55.805 ;
		RECT	0 56.105 0.32 56.805 ;
		RECT	0 57.105 0.32 57.595 ;
		RECT	0 57.895 0.32 58.08 ;
		RECT	0 58.38 0.32 58.485 ;
		RECT	0 58.785 0.32 59.25 ;
		RECT	0 59.55 0.32 59.625 ;
		RECT	0 59.925 0.32 60.08 ;
		RECT	0 60.58 0.32 61.825 ;
		RECT	0 62.125 0.32 62.25 ;
		RECT	0 62.76 0.32 63.14 ;
		RECT	0 63.44 0.32 65.28 ;
		RECT	0 65.58 0.32 65.685 ;
		RECT	0 65.985 0.32 66.17 ;
		RECT	0 66.725 0.32 67.2 ;
		RECT	0 67.5 0.32 69.81 ;
		RECT	0 70.11 0.32 70.205 ;
		RECT	0 70.505 0.32 70.75 ;
		RECT	0 71.05 0.32 72.365 ;
		RECT	0 72.925 0.32 73.355 ;
		RECT	0 73.655 0.32 75.245 ;
		RECT	0 75.805 0.32 76.235 ;
		RECT	0 76.535 0.32 78.125 ;
		RECT	0 78.685 0.32 79.115 ;
		RECT	0 79.415 0.32 81.005 ;
		RECT	0 81.565 0.32 81.995 ;
		RECT	0 82.295 0.32 83.885 ;
		RECT	0 84.445 0.32 84.875 ;
		RECT	0 85.175 0.32 86.765 ;
		RECT	0 87.325 0.32 87.755 ;
		RECT	0 88.055 0.32 89.645 ;
		RECT	0 90.205 0.32 90.635 ;
		RECT	0 90.935 0.32 92.525 ;
		RECT	0 93.085 0.32 93.515 ;
		RECT	0 93.815 0.32 95.405 ;
		RECT	0 95.965 0.32 96.395 ;
		RECT	0 96.695 0.32 98.285 ;
		RECT	0 98.845 0.32 99.275 ;
		RECT	0 99.575 0.32 100.38 ;
		RECT	20.845 0 21.165 100.94 ;
		RECT	0.32 0 20.845 0.35 ;
		RECT	0.32 100.59 20.845 100.94 ;
		LAYER	M3 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 20.845 100.59 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 1.665 0.32 2.095 ;
		RECT	0 2.655 0.32 4.245 ;
		RECT	0 4.545 0.32 4.975 ;
		RECT	0 5.535 0.32 7.125 ;
		RECT	0 7.425 0.32 7.855 ;
		RECT	0 8.415 0.32 10.005 ;
		RECT	0 10.305 0.32 10.735 ;
		RECT	0 11.295 0.32 12.885 ;
		RECT	0 13.185 0.32 13.615 ;
		RECT	0 14.175 0.32 15.765 ;
		RECT	0 16.065 0.32 16.495 ;
		RECT	0 17.055 0.32 18.645 ;
		RECT	0 18.945 0.32 19.375 ;
		RECT	0 19.935 0.32 21.525 ;
		RECT	0 21.825 0.32 22.255 ;
		RECT	0 22.815 0.32 24.405 ;
		RECT	0 24.705 0.32 25.135 ;
		RECT	0 25.695 0.32 28.6 ;
		RECT	0 28.9 0.32 28.95 ;
		RECT	0 29.25 0.32 29.61 ;
		RECT	0 30.31 0.32 31.95 ;
		RECT	0 32.555 0.32 32.77 ;
		RECT	0 33.07 0.32 33.175 ;
		RECT	0 33.475 0.32 35.285 ;
		RECT	0 35.585 0.32 35.8 ;
		RECT	0 36.1 0.32 36.205 ;
		RECT	0 36.505 0.32 38.345 ;
		RECT	0 38.645 0.32 38.83 ;
		RECT	0 39.13 0.32 39.235 ;
		RECT	0 39.535 0.32 39.63 ;
		RECT	0 39.93 0.32 40 ;
		RECT	0 40.3 0.32 40.375 ;
		RECT	0 40.675 0.32 40.86 ;
		RECT	0 41.57 0.32 43.005 ;
		RECT	0 43.705 0.32 43.89 ;
		RECT	0 44.475 0.32 47.4 ;
		RECT	0 48.1 0.32 48.57 ;
		RECT	0 48.87 0.32 50.235 ;
		RECT	0 50.535 0.32 54.325 ;
		RECT	0 54.86 0.32 55.05 ;
		RECT	0 55.35 0.32 55.425 ;
		RECT	0 55.725 0.32 55.805 ;
		RECT	0 56.105 0.32 56.805 ;
		RECT	0 57.105 0.32 57.595 ;
		RECT	0 57.895 0.32 58.08 ;
		RECT	0 58.38 0.32 58.485 ;
		RECT	0 58.785 0.32 59.25 ;
		RECT	0 59.55 0.32 59.625 ;
		RECT	0 59.925 0.32 60.08 ;
		RECT	0 60.58 0.32 61.825 ;
		RECT	0 62.125 0.32 62.25 ;
		RECT	0 62.76 0.32 63.14 ;
		RECT	0 63.44 0.32 65.28 ;
		RECT	0 65.58 0.32 65.685 ;
		RECT	0 65.985 0.32 66.17 ;
		RECT	0 66.725 0.32 67.2 ;
		RECT	0 67.5 0.32 69.81 ;
		RECT	0 70.11 0.32 70.205 ;
		RECT	0 70.505 0.32 70.75 ;
		RECT	0 71.05 0.32 72.365 ;
		RECT	0 72.925 0.32 73.355 ;
		RECT	0 73.655 0.32 75.245 ;
		RECT	0 75.805 0.32 76.235 ;
		RECT	0 76.535 0.32 78.125 ;
		RECT	0 78.685 0.32 79.115 ;
		RECT	0 79.415 0.32 81.005 ;
		RECT	0 81.565 0.32 81.995 ;
		RECT	0 82.295 0.32 83.885 ;
		RECT	0 84.445 0.32 84.875 ;
		RECT	0 85.175 0.32 86.765 ;
		RECT	0 87.325 0.32 87.755 ;
		RECT	0 88.055 0.32 89.645 ;
		RECT	0 90.205 0.32 90.635 ;
		RECT	0 90.935 0.32 92.525 ;
		RECT	0 93.085 0.32 93.515 ;
		RECT	0 93.815 0.32 95.405 ;
		RECT	0 95.965 0.32 96.395 ;
		RECT	0 96.695 0.32 98.285 ;
		RECT	0 98.845 0.32 99.275 ;
		RECT	0 99.575 0.32 100.38 ;
		RECT	20.845 0 21.165 100.94 ;
		RECT	0.32 0 20.845 0.35 ;
		RECT	0.32 100.59 20.845 100.94 ;
		LAYER	M4 DESIGNRULEWIDTH 0.165 ;
		RECT	0.57 26.775 14.49 27.945 ;
		RECT	14.185 27.945 14.49 28.175 ;
		RECT	0.57 28.005 14.125 28.155 ;
		RECT	0.57 28.905 14.49 29.015 ;
		RECT	0.57 29.15 14.49 29.34 ;
		RECT	0.57 29.825 14.49 29.925 ;
		RECT	0.57 30.315 11.56 30.415 ;
		RECT	0.57 30.805 14.49 30.905 ;
		RECT	11.255 30.905 14.49 30.91 ;
		RECT	11.255 30.91 12.345 31.255 ;
		RECT	0.57 31.005 11.155 31.215 ;
		RECT	12.445 31.01 14.49 31.2 ;
		RECT	11.255 31.255 11.56 31.315 ;
		RECT	0.57 31.315 11.56 31.385 ;
		RECT	0.57 31.485 14.49 31.675 ;
		RECT	0.57 31.775 14.49 31.93 ;
		RECT	0.57 32.32 14.49 32.385 ;
		RECT	0.57 32.775 14.49 32.88 ;
		RECT	0.57 33.27 14.49 33.37 ;
		RECT	0.57 33.76 14.15 33.86 ;
		RECT	0.57 34.25 14.49 34.355 ;
		RECT	0.57 34.745 14.49 34.845 ;
		RECT	0.57 35.235 14.49 35.34 ;
		RECT	0.57 35.44 14.49 35.63 ;
		RECT	0.57 35.73 14.49 35.83 ;
		RECT	0.57 36.22 14.49 36.325 ;
		RECT	0.57 36.715 14.49 36.815 ;
		RECT	0.57 37.205 14.49 37.305 ;
		RECT	0.57 37.695 14.49 37.8 ;
		RECT	0.57 38.19 14.49 38.29 ;
		RECT	0.57 38.68 14.49 38.78 ;
		RECT	0.57 39.17 14.49 39.275 ;
		RECT	0.57 39.375 14.49 39.565 ;
		RECT	0.57 39.665 14.49 39.765 ;
		RECT	0.57 40.155 14.49 40.26 ;
		RECT	0.57 40.65 14.49 40.75 ;
		RECT	8.61 41.14 14.49 41.23 ;
		RECT	0.57 41.155 8.56 41.225 ;
		RECT	0.57 41.64 14.49 41.735 ;
		RECT	0.57 42.125 14.49 42.225 ;
		RECT	0.57 42.615 14.49 42.72 ;
		RECT	9.515 43.11 14.49 43.2 ;
		RECT	9.295 43.115 9.465 43.125 ;
		RECT	0.57 43.125 9.465 43.195 ;
		RECT	9.295 43.195 9.465 43.205 ;
		RECT	0.57 43.3 14.49 43.51 ;
		RECT	0.57 43.61 14.49 43.705 ;
		RECT	0.57 44.095 14.49 44.2 ;
		RECT	0.57 44.59 14.49 44.685 ;
		RECT	0.57 45.075 14.49 45.18 ;
		RECT	0.57 45.57 14.49 45.655 ;
		RECT	0.57 46.045 14.49 46.28 ;
		RECT	0.57 46.28 13.465 46.395 ;
		RECT	13.565 46.38 14.49 46.57 ;
		RECT	11.215 46.395 13.465 46.655 ;
		RECT	0.57 46.455 11.155 46.605 ;
		RECT	0.57 47.045 13.8 47.145 ;
		RECT	0.57 47.245 14.49 47.435 ;
		RECT	0.57 47.535 13.8 47.64 ;
		RECT	0.57 48.03 14.49 48.13 ;
		RECT	0.57 48.52 14.49 48.62 ;
		RECT	0.57 49.01 7.02 49.115 ;
		RECT	13.595 49.01 14.49 49.115 ;
		RECT	0.57 49.505 14.49 49.605 ;
		RECT	0.57 49.995 14.49 50.1 ;
		RECT	0.57 50.49 13.8 50.59 ;
		RECT	0.57 50.69 14.49 50.88 ;
		RECT	0.57 50.98 13.8 51.08 ;
		RECT	11.215 51.47 13.5 51.73 ;
		RECT	13.6 51.495 14.49 51.685 ;
		RECT	0.57 51.52 11.155 51.67 ;
		RECT	0.57 51.73 13.5 51.785 ;
		RECT	0.57 51.785 14.49 52.08 ;
		RECT	0.57 52.47 14.49 52.555 ;
		RECT	0.57 52.945 14.49 53.05 ;
		RECT	0.57 53.44 14.49 53.545 ;
		RECT	0.57 53.935 14.49 54.025 ;
		RECT	7.785 54.435 14.49 54.515 ;
		RECT	0.57 54.44 7.735 54.51 ;
		RECT	0.57 54.615 14.49 54.825 ;
		RECT	0.57 54.925 14.49 55.02 ;
		RECT	0.57 55.41 14.49 55.51 ;
		RECT	0.57 55.9 14.49 56.005 ;
		RECT	0.57 56.395 14.49 56.485 ;
		RECT	8.06 56.895 14.49 56.985 ;
		RECT	0.57 56.9 8.01 56.97 ;
		RECT	0.57 57.375 14.49 57.48 ;
		RECT	0.57 57.87 14.49 57.97 ;
		RECT	0.57 58.36 14.49 58.465 ;
		RECT	0.57 58.565 14.49 58.755 ;
		RECT	0.57 58.855 14.49 58.955 ;
		RECT	0.57 59.345 14.49 59.445 ;
		RECT	0.57 59.835 14.49 59.94 ;
		RECT	0.57 60.33 14.49 60.43 ;
		RECT	0.57 60.82 14.49 60.925 ;
		RECT	0.57 61.315 14.49 61.415 ;
		RECT	0.57 61.805 14.49 61.905 ;
		RECT	0.57 62.295 14.15 62.39 ;
		RECT	0.57 62.49 14.49 62.7 ;
		RECT	2.785 62.8 14.49 62.89 ;
		RECT	0.57 63.28 14.49 63.375 ;
		RECT	0.57 63.79 14.49 63.86 ;
		RECT	0.57 64.28 14.49 64.35 ;
		RECT	0.57 64.765 14.49 64.825 ;
		RECT	0.57 65.215 14.49 65.35 ;
		RECT	0.57 65.74 14.49 65.81 ;
		RECT	0.57 66.2 14.49 66.35 ;
		RECT	0.57 66.45 14.49 66.64 ;
		RECT	0.57 66.74 12.555 66.815 ;
		RECT	11.255 66.815 12.555 66.825 ;
		RECT	11.255 66.825 12.27 67.215 ;
		RECT	0.57 66.915 11.155 67.125 ;
		RECT	12.37 66.925 14.49 67.115 ;
		RECT	11.255 67.215 14.49 67.225 ;
		RECT	0.57 67.225 14.49 67.32 ;
		RECT	0.57 67.71 12.555 67.81 ;
		RECT	0.57 68.2 14.49 68.305 ;
		RECT	0.57 68.705 14.49 68.915 ;
		RECT	0.57 69.045 14.49 69.155 ;
		RECT	14.21 69.885 14.49 70.115 ;
		RECT	0.57 69.905 14.15 70.055 ;
		RECT	0.57 70.115 14.49 71.285 ;
		RECT	0.21 28.005 0.57 28.155 ;
		RECT	0.215 29.15 0.57 29.34 ;
		RECT	0.22 31.005 0.57 31.215 ;
		RECT	0.22 31.485 0.57 31.675 ;
		RECT	0.22 35.44 0.57 35.63 ;
		RECT	0.23 39.375 0.57 39.565 ;
		RECT	0.14 41.155 0.57 41.225 ;
		RECT	0.15 43.125 0.57 43.195 ;
		RECT	0.215 43.3 0.57 43.51 ;
		RECT	0.21 46.455 0.57 46.605 ;
		RECT	0.225 47.245 0.57 47.435 ;
		RECT	0.325 50.69 0.61 50.88 ;
		RECT	0.21 51.52 0.57 51.67 ;
		RECT	0.15 54.44 0.57 54.51 ;
		RECT	0.235 54.615 0.57 54.825 ;
		RECT	0.14 56.9 0.57 56.97 ;
		RECT	0.24 58.565 0.57 58.755 ;
		RECT	0.225 62.49 0.57 62.7 ;
		RECT	0.14 62.805 0.57 62.875 ;
		RECT	0.235 66.45 0.57 66.64 ;
		RECT	0.225 66.915 0.57 67.125 ;
		RECT	0.24 68.705 0.57 68.915 ;
		RECT	0.22 69.905 0.57 70.055 ;
		RECT	5.7 23.225 13.945 23.375 ;
		RECT	5.7 20.345 13.945 20.495 ;
		RECT	5.7 17.465 13.945 17.615 ;
		RECT	5.7 14.585 13.945 14.735 ;
		RECT	5.7 11.705 13.945 11.855 ;
		RECT	5.7 8.825 13.945 8.975 ;
		RECT	5.7 5.945 13.945 6.095 ;
		RECT	5.7 3.065 13.945 3.215 ;
		RECT	5.7 26.105 13.945 26.255 ;
		RECT	0.57 23.225 1.11 23.375 ;
		RECT	0.57 20.345 1.11 20.495 ;
		RECT	0.57 17.465 1.11 17.615 ;
		RECT	0.57 14.585 1.11 14.735 ;
		RECT	0.57 11.705 1.11 11.855 ;
		RECT	0.57 8.825 1.11 8.975 ;
		RECT	0.57 5.945 1.11 6.095 ;
		RECT	0.57 3.065 1.11 3.215 ;
		RECT	0.57 26.105 1.11 26.255 ;
		RECT	1.005 23.225 5.7 23.375 ;
		RECT	1.005 20.345 5.7 20.495 ;
		RECT	1.005 17.465 5.7 17.615 ;
		RECT	1.005 14.585 5.7 14.735 ;
		RECT	1.005 11.705 5.7 11.855 ;
		RECT	1.005 8.825 5.7 8.975 ;
		RECT	1.005 5.945 5.7 6.095 ;
		RECT	1.005 3.065 5.7 3.215 ;
		RECT	1.005 26.105 5.7 26.255 ;
		RECT	0.255 26.105 0.57 26.255 ;
		RECT	0.255 23.225 0.57 23.375 ;
		RECT	0.255 20.345 0.57 20.495 ;
		RECT	0.255 17.465 0.57 17.615 ;
		RECT	0.255 14.585 0.57 14.735 ;
		RECT	0.255 11.705 0.57 11.855 ;
		RECT	0.255 8.825 0.57 8.975 ;
		RECT	0.255 5.945 0.57 6.095 ;
		RECT	0.255 3.065 0.57 3.215 ;
		RECT	5.7 74.685 13.945 74.835 ;
		RECT	5.7 77.565 13.945 77.715 ;
		RECT	5.7 80.445 13.945 80.595 ;
		RECT	5.7 83.325 13.945 83.475 ;
		RECT	5.7 86.205 13.945 86.355 ;
		RECT	5.7 89.085 13.945 89.235 ;
		RECT	5.7 91.965 13.945 92.115 ;
		RECT	5.7 94.845 13.945 94.995 ;
		RECT	5.7 97.725 13.945 97.875 ;
		RECT	5.7 71.805 13.945 71.955 ;
		RECT	0.57 74.685 1.11 74.835 ;
		RECT	0.57 77.565 1.11 77.715 ;
		RECT	0.57 80.445 1.11 80.595 ;
		RECT	0.57 83.325 1.11 83.475 ;
		RECT	0.57 86.205 1.11 86.355 ;
		RECT	0.57 89.085 1.11 89.235 ;
		RECT	0.57 91.965 1.11 92.115 ;
		RECT	0.57 94.845 1.11 94.995 ;
		RECT	0.57 97.725 1.11 97.875 ;
		RECT	0.57 71.805 1.11 71.955 ;
		RECT	1.005 74.685 5.7 74.835 ;
		RECT	1.005 77.565 5.7 77.715 ;
		RECT	1.005 80.445 5.7 80.595 ;
		RECT	1.005 83.325 5.7 83.475 ;
		RECT	1.005 86.205 5.7 86.355 ;
		RECT	1.005 89.085 5.7 89.235 ;
		RECT	1.005 91.965 5.7 92.115 ;
		RECT	1.005 94.845 5.7 94.995 ;
		RECT	1.005 97.725 5.7 97.875 ;
		RECT	1.005 71.805 5.7 71.955 ;
		RECT	0.255 71.805 0.57 71.955 ;
		RECT	0.255 74.685 0.57 74.835 ;
		RECT	0.255 77.565 0.57 77.715 ;
		RECT	0.255 80.445 0.57 80.595 ;
		RECT	0.255 83.325 0.57 83.475 ;
		RECT	0.255 86.205 0.57 86.355 ;
		RECT	0.255 89.085 0.57 89.235 ;
		RECT	0.255 91.965 0.57 92.115 ;
		RECT	0.255 94.845 0.57 94.995 ;
		RECT	0.255 97.725 0.57 97.875 ;
		RECT	15.63 28.905 16.17 29.015 ;
		RECT	15.63 26.775 16.17 28.175 ;
		RECT	16.17 28.905 16.71 29.015 ;
		RECT	16.17 26.775 16.71 28.175 ;
		RECT	16.71 28.905 17.25 29.015 ;
		RECT	16.71 26.775 17.25 28.175 ;
		RECT	15.09 28.905 15.63 29.015 ;
		RECT	15.09 26.775 15.63 28.175 ;
		RECT	14.49 28.905 15.09 29.015 ;
		RECT	14.49 26.775 15.09 28.175 ;
		RECT	17.25 28.905 17.79 29.015 ;
		RECT	17.25 26.775 17.79 28.175 ;
		RECT	17.79 28.905 18.33 29.015 ;
		RECT	17.79 26.775 18.33 28.175 ;
		RECT	18.33 28.905 18.87 29.015 ;
		RECT	18.33 26.775 18.87 28.175 ;
		RECT	19.41 28.905 20.01 29.015 ;
		RECT	19.41 26.775 20.01 28.175 ;
		RECT	18.87 28.905 19.41 29.015 ;
		RECT	18.87 26.775 19.41 28.175 ;
		RECT	15.09 69.045 15.63 69.155 ;
		RECT	15.09 69.885 15.63 71.285 ;
		RECT	14.49 69.045 15.09 69.155 ;
		RECT	14.49 69.885 15.09 71.285 ;
		RECT	15.63 69.045 16.17 69.155 ;
		RECT	15.63 69.885 16.17 71.285 ;
		RECT	16.17 69.045 16.71 69.155 ;
		RECT	16.17 69.885 16.71 71.285 ;
		RECT	16.71 69.045 17.25 69.155 ;
		RECT	16.71 69.885 17.25 71.285 ;
		RECT	17.25 69.045 17.79 69.155 ;
		RECT	17.25 69.885 17.79 71.285 ;
		RECT	17.79 69.045 18.33 69.155 ;
		RECT	17.79 69.885 18.33 71.285 ;
		RECT	18.33 69.045 18.87 69.155 ;
		RECT	18.33 69.885 18.87 71.285 ;
		RECT	19.41 69.045 20.01 69.155 ;
		RECT	19.41 69.885 20.01 71.285 ;
		RECT	18.87 69.045 19.41 69.155 ;
		RECT	18.87 69.885 19.41 71.285 ;
		RECT	20.01 26.775 21.165 28.175 ;
		RECT	20.01 28.905 21.165 29.015 ;
		RECT	20.97 29.015 21.165 29.435 ;
		RECT	20.01 29.15 20.87 29.34 ;
		RECT	20.01 29.825 21.165 29.925 ;
		RECT	20.01 30.805 21.165 30.91 ;
		RECT	20.97 30.91 21.165 31.255 ;
		RECT	20.01 31.01 20.87 31.2 ;
		RECT	20.97 31.435 21.165 31.775 ;
		RECT	20.01 31.485 20.87 31.675 ;
		RECT	20.92 31.775 21.165 31.93 ;
		RECT	20.01 31.78 20.86 31.93 ;
		RECT	20.01 32.32 21.165 32.385 ;
		RECT	20.01 32.775 21.165 32.88 ;
		RECT	20.01 33.27 21.165 33.37 ;
		RECT	20.41 33.76 21.165 33.86 ;
		RECT	20.01 34.25 21.165 34.355 ;
		RECT	20.79 34.355 21.165 34.745 ;
		RECT	20.01 34.745 21.165 34.845 ;
		RECT	20.01 35.235 21.165 35.34 ;
		RECT	20.97 35.34 21.165 35.73 ;
		RECT	20.01 35.44 20.87 35.63 ;
		RECT	20.01 35.73 21.165 35.83 ;
		RECT	20.01 36.22 21.165 36.325 ;
		RECT	20.01 36.715 21.165 36.815 ;
		RECT	20.01 37.205 21.165 37.305 ;
		RECT	20.01 37.695 21.165 37.8 ;
		RECT	20.01 38.19 21.165 38.29 ;
		RECT	20.01 38.68 21.165 38.78 ;
		RECT	20.01 39.17 21.165 39.275 ;
		RECT	20.97 39.275 21.165 39.665 ;
		RECT	20.01 39.375 20.87 39.565 ;
		RECT	20.01 39.665 21.165 39.765 ;
		RECT	20.01 40.155 21.165 40.26 ;
		RECT	20.01 40.65 21.165 40.75 ;
		RECT	20.01 41.14 21.165 41.23 ;
		RECT	20.01 41.64 21.165 41.735 ;
		RECT	20.01 42.125 21.165 42.225 ;
		RECT	20.01 42.615 21.165 42.72 ;
		RECT	20.01 43.11 21.165 43.2 ;
		RECT	20.97 43.2 21.165 43.61 ;
		RECT	20.01 43.3 20.87 43.51 ;
		RECT	20.01 43.61 21.165 43.705 ;
		RECT	20.97 43.705 21.165 44.095 ;
		RECT	20.01 44.095 21.165 44.2 ;
		RECT	20.01 44.59 21.165 44.685 ;
		RECT	20.01 45.075 21.165 45.18 ;
		RECT	20.01 45.57 21.165 45.655 ;
		RECT	20.97 45.655 21.165 46.655 ;
		RECT	20.01 46.055 20.87 46.265 ;
		RECT	20.01 46.38 20.86 46.57 ;
		RECT	20.97 47.19 21.165 47.495 ;
		RECT	20.01 47.245 20.87 47.435 ;
		RECT	20.01 48.03 21.165 48.13 ;
		RECT	20.01 48.52 21.165 48.62 ;
		RECT	20.01 49.01 21.165 49.115 ;
		RECT	20.01 49.505 21.165 49.605 ;
		RECT	20.01 49.995 21.165 50.1 ;
		RECT	20.97 50.635 21.165 50.935 ;
		RECT	20.01 50.69 20.87 50.88 ;
		RECT	20.97 51.47 21.165 52.47 ;
		RECT	20.01 51.495 20.87 51.685 ;
		RECT	20.01 51.83 20.87 52.04 ;
		RECT	20.01 52.47 21.165 52.555 ;
		RECT	20.01 52.945 21.165 53.05 ;
		RECT	20.01 53.44 21.165 53.545 ;
		RECT	20.01 53.935 21.165 54.025 ;
		RECT	20.97 54.025 21.165 54.435 ;
		RECT	20.01 54.435 21.165 54.515 ;
		RECT	20.97 54.515 21.165 54.925 ;
		RECT	20.01 54.615 20.87 54.825 ;
		RECT	20.01 54.925 21.165 55.02 ;
		RECT	20.01 55.41 21.165 55.51 ;
		RECT	20.01 55.9 21.165 56.005 ;
		RECT	20.01 56.395 21.165 56.485 ;
		RECT	20.01 56.895 21.165 56.985 ;
		RECT	20.01 57.375 21.165 57.48 ;
		RECT	20.01 57.87 21.165 57.97 ;
		RECT	20.01 58.36 21.165 58.465 ;
		RECT	20.97 58.465 21.165 58.855 ;
		RECT	20.01 58.565 20.87 58.755 ;
		RECT	20.01 58.855 21.165 58.955 ;
		RECT	20.01 59.345 21.165 59.445 ;
		RECT	20.01 59.835 21.165 59.94 ;
		RECT	20.01 60.33 21.165 60.43 ;
		RECT	20.01 60.82 21.165 60.925 ;
		RECT	20.01 61.315 21.165 61.415 ;
		RECT	20.01 61.805 21.165 61.905 ;
		RECT	20.41 62.295 21.165 62.39 ;
		RECT	20.97 62.39 21.165 62.8 ;
		RECT	20.01 62.49 20.87 62.7 ;
		RECT	20.01 62.8 21.165 62.89 ;
		RECT	20.01 63.28 21.165 63.375 ;
		RECT	20.79 63.375 21.165 63.785 ;
		RECT	20.74 63.785 21.165 63.875 ;
		RECT	20.74 64.265 21.165 64.355 ;
		RECT	20.01 64.765 21.165 64.825 ;
		RECT	20.01 65.215 21.165 65.35 ;
		RECT	20.01 65.74 21.165 65.81 ;
		RECT	20.97 66.2 21.165 66.69 ;
		RECT	20.01 66.2 20.87 66.35 ;
		RECT	20.01 66.45 20.87 66.64 ;
		RECT	20.97 66.87 21.165 67.215 ;
		RECT	20.01 66.925 20.87 67.115 ;
		RECT	20.01 67.215 21.165 67.32 ;
		RECT	20.01 68.2 21.165 68.305 ;
		RECT	20.97 68.695 21.165 69.045 ;
		RECT	20.01 68.705 20.87 68.915 ;
		RECT	20.01 69.045 21.165 69.155 ;
		RECT	20.01 69.885 21.165 71.285 ;
		RECT	14.49 29.15 19.41 29.34 ;
		RECT	14.49 29.825 19.41 29.925 ;
		RECT	14.49 30.805 19.41 30.91 ;
		RECT	14.49 31.01 19.41 31.2 ;
		RECT	14.49 31.485 19.41 31.675 ;
		RECT	14.59 31.78 19.41 31.93 ;
		RECT	14.49 32.32 19.41 32.385 ;
		RECT	14.49 32.775 19.41 32.88 ;
		RECT	14.49 33.27 19.41 33.37 ;
		RECT	14.49 34.25 19.41 34.355 ;
		RECT	14.49 34.745 19.41 34.845 ;
		RECT	14.49 35.235 19.41 35.34 ;
		RECT	14.49 35.44 19.41 35.63 ;
		RECT	14.49 35.73 19.41 35.83 ;
		RECT	14.49 36.22 19.41 36.325 ;
		RECT	14.49 36.715 19.41 36.815 ;
		RECT	14.49 37.205 19.41 37.305 ;
		RECT	14.49 37.695 19.41 37.8 ;
		RECT	14.49 38.19 19.41 38.29 ;
		RECT	14.49 38.68 19.41 38.78 ;
		RECT	14.49 39.17 19.41 39.275 ;
		RECT	14.49 39.375 19.41 39.565 ;
		RECT	14.49 39.665 19.41 39.765 ;
		RECT	14.49 40.155 19.41 40.26 ;
		RECT	14.49 40.65 19.41 40.75 ;
		RECT	14.49 41.14 19.41 41.23 ;
		RECT	14.49 41.64 19.41 41.735 ;
		RECT	14.49 42.125 19.41 42.225 ;
		RECT	14.49 42.615 19.41 42.72 ;
		RECT	14.49 43.11 19.41 43.2 ;
		RECT	14.49 43.3 19.41 43.51 ;
		RECT	14.49 43.61 19.41 43.705 ;
		RECT	14.49 44.095 19.41 44.2 ;
		RECT	14.49 44.59 19.41 44.685 ;
		RECT	14.49 45.075 19.41 45.18 ;
		RECT	14.49 45.57 19.41 45.655 ;
		RECT	14.49 46.045 14.595 46.28 ;
		RECT	14.695 46.055 19.41 46.265 ;
		RECT	14.49 46.38 19.41 46.57 ;
		RECT	14.49 47.245 19.41 47.435 ;
		RECT	14.49 48.03 19.41 48.13 ;
		RECT	14.49 48.52 19.41 48.62 ;
		RECT	14.49 49.01 19.41 49.115 ;
		RECT	14.49 49.505 19.41 49.605 ;
		RECT	14.49 49.995 19.41 50.1 ;
		RECT	14.49 50.69 19.41 50.88 ;
		RECT	14.49 51.495 19.41 51.685 ;
		RECT	14.59 51.83 19.41 52.04 ;
		RECT	14.49 52.47 19.41 52.555 ;
		RECT	14.49 52.945 19.41 53.05 ;
		RECT	14.49 53.44 19.41 53.545 ;
		RECT	14.49 53.935 19.41 54.025 ;
		RECT	14.49 54.435 19.41 54.515 ;
		RECT	14.49 54.615 19.41 54.825 ;
		RECT	14.49 54.925 19.41 55.02 ;
		RECT	14.49 55.41 19.41 55.51 ;
		RECT	14.49 55.9 19.41 56.005 ;
		RECT	14.49 56.395 19.41 56.485 ;
		RECT	14.49 56.895 19.41 56.985 ;
		RECT	14.49 57.375 19.41 57.48 ;
		RECT	14.49 57.87 19.41 57.97 ;
		RECT	14.49 58.36 19.41 58.465 ;
		RECT	14.49 58.565 19.41 58.755 ;
		RECT	14.49 58.855 19.41 58.955 ;
		RECT	14.49 59.345 19.41 59.445 ;
		RECT	14.49 59.835 19.41 59.94 ;
		RECT	14.49 60.33 19.41 60.43 ;
		RECT	14.49 60.82 19.41 60.925 ;
		RECT	14.49 61.315 19.41 61.415 ;
		RECT	14.49 61.805 19.41 61.905 ;
		RECT	14.49 62.49 19.41 62.7 ;
		RECT	14.49 62.8 19.41 62.89 ;
		RECT	14.49 63.28 19.41 63.375 ;
		RECT	14.49 63.79 19.41 63.86 ;
		RECT	14.49 64.28 19.445 64.35 ;
		RECT	14.49 64.765 19.41 64.825 ;
		RECT	14.49 65.215 19.41 65.35 ;
		RECT	14.49 65.74 19.41 65.81 ;
		RECT	14.49 66.2 14.63 66.35 ;
		RECT	14.69 66.2 19.41 66.35 ;
		RECT	14.49 66.45 19.41 66.64 ;
		RECT	14.49 66.925 19.41 67.115 ;
		RECT	14.49 67.215 19.41 67.32 ;
		RECT	14.49 68.2 19.41 68.305 ;
		RECT	14.49 68.705 19.41 68.915 ;
		RECT	19.41 29.15 20.01 29.34 ;
		RECT	19.41 29.825 20.01 29.925 ;
		RECT	19.41 30.805 20.01 30.91 ;
		RECT	19.41 31.01 20.01 31.2 ;
		RECT	19.41 31.485 20.01 31.675 ;
		RECT	19.41 31.78 20.175 31.93 ;
		RECT	19.41 32.32 20.01 32.385 ;
		RECT	19.41 32.775 20.01 32.88 ;
		RECT	19.41 33.27 20.01 33.37 ;
		RECT	19.41 34.25 20.01 34.355 ;
		RECT	19.41 34.745 20.01 34.845 ;
		RECT	19.41 35.235 20.01 35.34 ;
		RECT	19.41 35.44 20.01 35.63 ;
		RECT	19.41 35.73 20.01 35.83 ;
		RECT	19.41 36.22 20.01 36.325 ;
		RECT	19.41 36.715 20.01 36.815 ;
		RECT	19.41 37.205 20.01 37.305 ;
		RECT	19.41 37.695 20.01 37.8 ;
		RECT	19.41 38.19 20.01 38.29 ;
		RECT	19.41 38.68 20.01 38.78 ;
		RECT	19.41 39.17 20.01 39.275 ;
		RECT	19.41 39.375 20.01 39.565 ;
		RECT	19.41 39.665 20.01 39.765 ;
		RECT	19.41 40.155 20.01 40.26 ;
		RECT	19.41 40.65 20.01 40.75 ;
		RECT	19.41 41.14 20.01 41.23 ;
		RECT	19.41 41.64 20.01 41.735 ;
		RECT	19.41 42.125 20.01 42.225 ;
		RECT	19.41 42.615 20.01 42.72 ;
		RECT	19.41 43.11 20.01 43.2 ;
		RECT	19.41 43.3 20.01 43.51 ;
		RECT	19.41 43.61 20.01 43.705 ;
		RECT	19.41 44.095 20.01 44.2 ;
		RECT	19.41 44.59 20.01 44.685 ;
		RECT	19.41 45.075 20.01 45.18 ;
		RECT	19.41 45.57 20.01 45.655 ;
		RECT	19.41 46.055 20.085 46.265 ;
		RECT	19.41 46.38 20.01 46.57 ;
		RECT	19.41 47.245 20.01 47.435 ;
		RECT	19.41 48.03 20.01 48.13 ;
		RECT	19.41 48.52 20.01 48.62 ;
		RECT	19.41 49.01 20.01 49.115 ;
		RECT	19.41 49.505 20.01 49.605 ;
		RECT	19.41 49.995 20.01 50.1 ;
		RECT	19.41 50.69 20.01 50.88 ;
		RECT	19.41 51.495 20.01 51.685 ;
		RECT	19.41 51.83 20.01 52.04 ;
		RECT	19.41 52.47 20.01 52.555 ;
		RECT	19.41 52.945 20.01 53.05 ;
		RECT	19.41 53.44 20.01 53.545 ;
		RECT	19.41 53.935 20.01 54.025 ;
		RECT	19.41 54.435 20.01 54.515 ;
		RECT	19.41 54.615 20.01 54.825 ;
		RECT	19.41 54.925 20.01 55.02 ;
		RECT	19.41 55.41 20.01 55.51 ;
		RECT	19.41 55.9 20.01 56.005 ;
		RECT	19.41 56.395 20.01 56.485 ;
		RECT	19.41 56.895 20.01 56.985 ;
		RECT	19.41 57.375 20.01 57.48 ;
		RECT	19.41 57.87 20.01 57.97 ;
		RECT	19.41 58.36 20.01 58.465 ;
		RECT	19.41 58.565 20.01 58.755 ;
		RECT	19.41 58.855 20.01 58.955 ;
		RECT	19.41 59.345 20.01 59.445 ;
		RECT	19.41 59.835 20.01 59.94 ;
		RECT	19.41 60.33 20.01 60.43 ;
		RECT	19.41 60.82 20.01 60.925 ;
		RECT	19.41 61.315 20.01 61.415 ;
		RECT	19.41 61.805 20.01 61.905 ;
		RECT	19.41 62.49 20.01 62.7 ;
		RECT	19.41 62.8 20.01 62.89 ;
		RECT	19.41 63.28 20.01 63.375 ;
		RECT	19.41 63.79 20.01 63.86 ;
		RECT	19.41 64.28 20.01 64.35 ;
		RECT	19.41 64.765 20.01 64.825 ;
		RECT	19.41 65.215 20.01 65.35 ;
		RECT	19.41 65.74 20.01 65.81 ;
		RECT	19.41 66.2 20.01 66.35 ;
		RECT	19.41 66.45 20.01 66.64 ;
		RECT	19.41 66.925 20.01 67.115 ;
		RECT	19.41 67.215 20.01 67.32 ;
		RECT	19.41 68.2 20.01 68.305 ;
		RECT	19.41 68.705 20.01 68.915 ;
		RECT	0.295 34.455 20.69 34.645 ;
		RECT	0.215 43.805 20.87 43.995 ;
		RECT	0.21 45.755 20.86 45.945 ;
		RECT	0.22 52.18 20.87 52.37 ;
		RECT	0.225 54.125 20.87 54.335 ;
		RECT	0.225 63.475 20.69 63.685 ;
		RECT	0.225 63.79 0.57 63.86 ;
		RECT	0.22 64.28 0.57 64.35 ;
		RECT	11.61 30.32 21.07 30.41 ;
		RECT	11.61 31.305 21.07 31.385 ;
		RECT	14.2 33.765 20.36 33.855 ;
		RECT	13.85 47.05 21.07 47.14 ;
		RECT	13.85 47.545 21.07 47.635 ;
		RECT	7.07 49.015 13.545 49.115 ;
		RECT	13.85 50.495 21.07 50.585 ;
		RECT	13.85 50.985 21.07 51.075 ;
		RECT	14.2 62.3 20.36 62.39 ;
		RECT	0.57 62.805 2.735 62.875 ;
		RECT	12.605 66.74 21.07 66.82 ;
		RECT	12.605 67.715 21.07 67.805 ;
		RECT	20.01 63.79 20.69 63.86 ;
		RECT	20.01 64.28 20.69 64.35 ;
		LAYER	VIA1 DESIGNRULEWIDTH 0.07 ;
		RECT	0 0 21.165 100.94 ;
		LAYER	VIA2 DESIGNRULEWIDTH 0.07 ;
		RECT	0 0 21.165 100.94 ;
		LAYER	VIA3 DESIGNRULEWIDTH 0.07 ;
		RECT	0.435 28.015 0.485 28.145 ;
		RECT	0.435 29.18 0.485 29.31 ;
		RECT	0.435 31.045 0.485 31.175 ;
		RECT	0.435 31.515 0.485 31.645 ;
		RECT	0.435 35.47 0.485 35.6 ;
		RECT	0.435 39.405 0.485 39.535 ;
		RECT	0.435 43.34 0.485 43.47 ;
		RECT	0.435 46.465 0.485 46.595 ;
		RECT	0.435 47.275 0.485 47.405 ;
		RECT	0.435 50.72 0.485 50.85 ;
		RECT	0.435 51.53 0.485 51.66 ;
		RECT	0.435 54.655 0.485 54.785 ;
		RECT	0.435 58.595 0.485 58.725 ;
		RECT	0.435 62.53 0.485 62.66 ;
		RECT	0.435 66.48 0.485 66.61 ;
		RECT	0.435 66.955 0.485 67.085 ;
		RECT	0.435 68.745 0.485 68.875 ;
		RECT	0.435 69.915 0.485 70.045 ;
		RECT	0.435 28.475 0.485 28.605 ;
		RECT	0.435 34.485 0.485 34.615 ;
		RECT	0.435 63.515 0.485 63.645 ;
		RECT	0.435 69.455 0.485 69.585 ;
		RECT	1.085 28.015 1.135 28.145 ;
		RECT	1.38 28.015 1.43 28.145 ;
		RECT	1.86 28.015 1.91 28.145 ;
		RECT	2.01 28.015 2.06 28.145 ;
		RECT	3.25 28.015 3.3 28.145 ;
		RECT	3.515 28.015 3.565 28.145 ;
		RECT	4.51 28.015 4.56 28.145 ;
		RECT	5.035 28.015 5.085 28.145 ;
		RECT	6.22 28.015 6.27 28.145 ;
		RECT	7.5 28.015 7.55 28.145 ;
		RECT	9.315 28.015 9.365 28.145 ;
		RECT	9.72 28.015 9.77 28.145 ;
		RECT	11.025 28.015 11.075 28.145 ;
		RECT	0.62 28.245 0.67 28.375 ;
		RECT	3.65 28.245 3.7 28.375 ;
		RECT	7.19 28.245 7.24 28.375 ;
		RECT	14.14 28.245 14.19 28.375 ;
		RECT	2.18 28.475 2.23 28.605 ;
		RECT	8.56 28.475 8.61 28.605 ;
		RECT	10.27 28.475 10.32 28.605 ;
		RECT	13.8 28.705 13.85 28.835 ;
		RECT	1.045 29.155 1.175 29.205 ;
		RECT	1.34 29.155 1.47 29.205 ;
		RECT	4.47 29.155 4.6 29.205 ;
		RECT	9.275 29.155 9.405 29.205 ;
		RECT	1.86 29.18 1.91 29.31 ;
		RECT	2.01 29.18 2.06 29.31 ;
		RECT	3.25 29.18 3.3 29.31 ;
		RECT	3.515 29.18 3.565 29.31 ;
		RECT	5.035 29.18 5.085 29.31 ;
		RECT	6.22 29.18 6.27 29.31 ;
		RECT	7.5 29.18 7.55 29.31 ;
		RECT	9.72 29.18 9.77 29.31 ;
		RECT	11.025 29.18 11.075 29.31 ;
		RECT	1.045 29.285 1.175 29.335 ;
		RECT	1.34 29.285 1.47 29.335 ;
		RECT	4.47 29.285 4.6 29.335 ;
		RECT	9.275 29.285 9.405 29.335 ;
		RECT	3.02 29.54 3.15 29.59 ;
		RECT	1.57 29.565 1.62 29.695 ;
		RECT	4.87 29.565 4.92 29.695 ;
		RECT	5.9 29.565 5.95 29.695 ;
		RECT	8.955 29.565 9.005 29.695 ;
		RECT	12.79 29.565 12.84 29.695 ;
		RECT	14.33 29.565 14.38 29.695 ;
		RECT	3.02 29.67 3.15 29.72 ;
		RECT	3.8 30.03 3.93 30.08 ;
		RECT	5.635 30.03 5.765 30.08 ;
		RECT	8.31 30.03 8.44 30.08 ;
		RECT	8.73 30.03 8.86 30.08 ;
		RECT	0.9 30.055 0.95 30.185 ;
		RECT	2.485 30.055 2.535 30.185 ;
		RECT	2.615 30.055 2.665 30.185 ;
		RECT	6.065 30.055 6.115 30.185 ;
		RECT	6.725 30.055 6.775 30.185 ;
		RECT	11.555 30.055 11.865 30.185 ;
		RECT	12.52 30.055 12.57 30.185 ;
		RECT	14.005 30.055 14.055 30.185 ;
		RECT	3.8 30.16 3.93 30.21 ;
		RECT	5.635 30.16 5.765 30.21 ;
		RECT	8.31 30.16 8.44 30.21 ;
		RECT	8.73 30.16 8.86 30.21 ;
		RECT	11.685 30.34 11.735 30.39 ;
		RECT	12.655 30.34 12.705 30.39 ;
		RECT	3.02 30.52 3.15 30.57 ;
		RECT	1.57 30.545 1.62 30.675 ;
		RECT	4.87 30.545 4.92 30.675 ;
		RECT	5.9 30.545 5.95 30.675 ;
		RECT	8.955 30.545 9.005 30.675 ;
		RECT	12.79 30.545 12.84 30.675 ;
		RECT	14.335 30.545 14.385 30.675 ;
		RECT	3.02 30.65 3.15 30.7 ;
		RECT	1.045 31.02 1.175 31.07 ;
		RECT	1.34 31.02 1.47 31.07 ;
		RECT	4.47 31.02 4.6 31.07 ;
		RECT	9.275 31.02 9.405 31.07 ;
		RECT	13.675 31.04 13.725 31.17 ;
		RECT	1.86 31.045 1.91 31.175 ;
		RECT	2.01 31.045 2.06 31.175 ;
		RECT	3.25 31.045 3.3 31.175 ;
		RECT	3.515 31.045 3.565 31.175 ;
		RECT	5.035 31.045 5.085 31.175 ;
		RECT	6.22 31.045 6.27 31.175 ;
		RECT	7.5 31.045 7.55 31.175 ;
		RECT	9.72 31.045 9.77 31.175 ;
		RECT	11.025 31.045 11.075 31.175 ;
		RECT	1.045 31.15 1.175 31.2 ;
		RECT	1.34 31.15 1.47 31.2 ;
		RECT	4.47 31.15 4.6 31.2 ;
		RECT	9.275 31.15 9.405 31.2 ;
		RECT	11.685 31.32 11.735 31.37 ;
		RECT	12.655 31.32 12.705 31.37 ;
		RECT	1.045 31.49 1.175 31.54 ;
		RECT	1.34 31.49 1.47 31.54 ;
		RECT	4.47 31.49 4.6 31.54 ;
		RECT	9.275 31.49 9.405 31.54 ;
		RECT	1.86 31.515 1.91 31.645 ;
		RECT	2.01 31.515 2.06 31.645 ;
		RECT	3.25 31.515 3.3 31.645 ;
		RECT	3.515 31.515 3.565 31.645 ;
		RECT	5.035 31.515 5.085 31.645 ;
		RECT	6.22 31.515 6.27 31.645 ;
		RECT	7.5 31.515 7.55 31.645 ;
		RECT	9.72 31.515 9.77 31.645 ;
		RECT	11.025 31.515 11.075 31.645 ;
		RECT	1.045 31.62 1.175 31.67 ;
		RECT	1.34 31.62 1.47 31.67 ;
		RECT	4.47 31.62 4.6 31.67 ;
		RECT	9.275 31.62 9.405 31.67 ;
		RECT	3.8 32.035 3.93 32.085 ;
		RECT	5.635 32.035 5.765 32.085 ;
		RECT	8.31 32.035 8.44 32.085 ;
		RECT	8.73 32.035 8.86 32.085 ;
		RECT	0.9 32.06 0.95 32.19 ;
		RECT	2.485 32.06 2.535 32.19 ;
		RECT	2.615 32.06 2.665 32.19 ;
		RECT	6.065 32.06 6.115 32.19 ;
		RECT	6.725 32.06 6.775 32.19 ;
		RECT	11.555 32.06 11.865 32.19 ;
		RECT	12.52 32.06 12.57 32.19 ;
		RECT	14.005 32.06 14.055 32.19 ;
		RECT	3.8 32.165 3.93 32.215 ;
		RECT	5.635 32.165 5.765 32.215 ;
		RECT	8.31 32.165 8.44 32.215 ;
		RECT	8.73 32.165 8.86 32.215 ;
		RECT	3.02 32.49 3.15 32.54 ;
		RECT	1.57 32.515 1.62 32.645 ;
		RECT	4.87 32.515 4.92 32.645 ;
		RECT	5.9 32.515 5.95 32.645 ;
		RECT	8.955 32.515 9.005 32.645 ;
		RECT	12.79 32.515 12.84 32.645 ;
		RECT	14.335 32.515 14.385 32.645 ;
		RECT	3.02 32.62 3.15 32.67 ;
		RECT	4.035 33.01 4.085 33.14 ;
		RECT	6.495 33.01 6.545 33.14 ;
		RECT	11.685 33.01 11.735 33.14 ;
		RECT	12.655 33.01 12.705 33.14 ;
		RECT	3.02 33.475 3.15 33.525 ;
		RECT	1.57 33.5 1.62 33.63 ;
		RECT	4.87 33.5 4.92 33.63 ;
		RECT	5.9 33.5 5.95 33.63 ;
		RECT	8.955 33.5 9.005 33.63 ;
		RECT	12.79 33.5 12.84 33.63 ;
		RECT	14.335 33.5 14.385 33.63 ;
		RECT	3.02 33.605 3.15 33.655 ;
		RECT	14.29 33.785 14.42 33.835 ;
		RECT	4.035 33.99 4.085 34.12 ;
		RECT	6.495 33.99 6.545 34.12 ;
		RECT	2.18 34.485 2.23 34.615 ;
		RECT	8.56 34.485 8.61 34.615 ;
		RECT	10.27 34.485 10.32 34.615 ;
		RECT	3.8 34.95 3.93 35 ;
		RECT	5.635 34.95 5.765 35 ;
		RECT	8.31 34.95 8.44 35 ;
		RECT	8.73 34.95 8.86 35 ;
		RECT	0.9 34.975 0.95 35.105 ;
		RECT	2.485 34.975 2.535 35.105 ;
		RECT	2.615 34.975 2.665 35.105 ;
		RECT	6.065 34.975 6.115 35.105 ;
		RECT	6.725 34.975 6.775 35.105 ;
		RECT	11.555 34.975 11.865 35.105 ;
		RECT	12.52 34.975 12.57 35.105 ;
		RECT	14.005 34.975 14.055 35.105 ;
		RECT	3.8 35.08 3.93 35.13 ;
		RECT	5.635 35.08 5.765 35.13 ;
		RECT	8.31 35.08 8.44 35.13 ;
		RECT	8.73 35.08 8.86 35.13 ;
		RECT	1.045 35.445 1.175 35.495 ;
		RECT	1.34 35.445 1.47 35.495 ;
		RECT	4.47 35.445 4.6 35.495 ;
		RECT	1.86 35.47 1.91 35.6 ;
		RECT	2.01 35.47 2.06 35.6 ;
		RECT	2.32 35.47 2.37 35.6 ;
		RECT	3.25 35.47 3.3 35.6 ;
		RECT	3.515 35.47 3.565 35.6 ;
		RECT	5.035 35.47 5.085 35.6 ;
		RECT	6.22 35.47 6.27 35.6 ;
		RECT	7.5 35.47 7.55 35.6 ;
		RECT	9.72 35.47 9.77 35.6 ;
		RECT	11.025 35.47 11.075 35.6 ;
		RECT	1.045 35.575 1.175 35.625 ;
		RECT	1.34 35.575 1.47 35.625 ;
		RECT	4.47 35.575 4.6 35.625 ;
		RECT	3.8 35.935 3.93 35.985 ;
		RECT	5.635 35.935 5.765 35.985 ;
		RECT	8.31 35.935 8.44 35.985 ;
		RECT	8.73 35.935 8.86 35.985 ;
		RECT	0.9 35.96 0.95 36.09 ;
		RECT	2.485 35.96 2.535 36.09 ;
		RECT	2.615 35.96 2.665 36.09 ;
		RECT	6.065 35.96 6.115 36.09 ;
		RECT	6.725 35.96 6.775 36.09 ;
		RECT	11.555 35.96 11.865 36.09 ;
		RECT	12.52 35.96 12.57 36.09 ;
		RECT	14.005 35.96 14.055 36.09 ;
		RECT	3.8 36.065 3.93 36.115 ;
		RECT	5.635 36.065 5.765 36.115 ;
		RECT	8.31 36.065 8.44 36.115 ;
		RECT	8.73 36.065 8.86 36.115 ;
		RECT	3.02 36.43 3.15 36.48 ;
		RECT	1.57 36.455 1.62 36.585 ;
		RECT	4.87 36.455 4.92 36.585 ;
		RECT	5.9 36.455 5.95 36.585 ;
		RECT	9.195 36.455 9.245 36.585 ;
		RECT	10.27 36.455 10.32 36.585 ;
		RECT	12.79 36.455 12.84 36.585 ;
		RECT	14.335 36.455 14.385 36.585 ;
		RECT	3.02 36.56 3.15 36.61 ;
		RECT	4.035 36.945 4.085 37.075 ;
		RECT	3.02 37.41 3.15 37.46 ;
		RECT	1.57 37.435 1.62 37.565 ;
		RECT	4.87 37.435 4.92 37.565 ;
		RECT	5.9 37.435 5.95 37.565 ;
		RECT	9.195 37.435 9.245 37.565 ;
		RECT	9.43 37.435 9.48 37.565 ;
		RECT	10.27 37.435 10.32 37.565 ;
		RECT	12.79 37.435 12.84 37.565 ;
		RECT	14.335 37.435 14.385 37.565 ;
		RECT	3.02 37.54 3.15 37.59 ;
		RECT	0.9 37.905 14.055 38.085 ;
		RECT	3.02 38.395 3.15 38.445 ;
		RECT	1.57 38.42 1.62 38.55 ;
		RECT	4.87 38.42 4.92 38.55 ;
		RECT	5.9 38.42 5.95 38.55 ;
		RECT	9.43 38.42 9.48 38.55 ;
		RECT	10.27 38.42 10.32 38.55 ;
		RECT	12.79 38.42 12.84 38.55 ;
		RECT	14.33 38.42 14.38 38.55 ;
		RECT	3.02 38.525 3.15 38.575 ;
		RECT	3.8 38.885 3.93 38.935 ;
		RECT	5.635 38.885 5.765 38.935 ;
		RECT	8.31 38.885 8.44 38.935 ;
		RECT	8.73 38.885 8.86 38.935 ;
		RECT	0.9 38.91 0.95 39.04 ;
		RECT	2.485 38.91 2.535 39.04 ;
		RECT	2.615 38.91 2.665 39.04 ;
		RECT	6.065 38.91 6.115 39.04 ;
		RECT	6.725 38.91 6.775 39.04 ;
		RECT	11.555 38.91 11.865 39.04 ;
		RECT	12.52 38.91 12.57 39.04 ;
		RECT	14.005 38.91 14.055 39.04 ;
		RECT	3.8 39.015 3.93 39.065 ;
		RECT	5.635 39.015 5.765 39.065 ;
		RECT	8.31 39.015 8.44 39.065 ;
		RECT	8.73 39.015 8.86 39.065 ;
		RECT	1.045 39.38 1.175 39.43 ;
		RECT	1.34 39.38 1.47 39.43 ;
		RECT	4.47 39.38 4.6 39.43 ;
		RECT	1.86 39.405 1.91 39.535 ;
		RECT	2.01 39.405 2.06 39.535 ;
		RECT	2.32 39.405 2.37 39.535 ;
		RECT	3.25 39.405 3.3 39.535 ;
		RECT	3.515 39.405 3.565 39.535 ;
		RECT	5.035 39.405 5.085 39.535 ;
		RECT	6.22 39.405 6.27 39.535 ;
		RECT	7.5 39.405 7.55 39.535 ;
		RECT	9.72 39.405 9.77 39.535 ;
		RECT	11.025 39.405 11.075 39.535 ;
		RECT	1.045 39.51 1.175 39.56 ;
		RECT	1.34 39.51 1.47 39.56 ;
		RECT	4.47 39.51 4.6 39.56 ;
		RECT	3.8 39.87 3.93 39.92 ;
		RECT	5.635 39.87 5.765 39.92 ;
		RECT	8.31 39.87 8.44 39.92 ;
		RECT	8.73 39.87 8.86 39.92 ;
		RECT	0.9 39.895 0.95 40.025 ;
		RECT	2.485 39.895 2.535 40.025 ;
		RECT	2.615 39.895 2.665 40.025 ;
		RECT	6.065 39.895 6.115 40.025 ;
		RECT	6.725 39.895 6.775 40.025 ;
		RECT	11.555 39.895 11.865 40.025 ;
		RECT	12.52 39.895 12.57 40.025 ;
		RECT	14.005 39.895 14.055 40.025 ;
		RECT	3.8 40 3.93 40.05 ;
		RECT	5.635 40 5.765 40.05 ;
		RECT	8.31 40 8.44 40.05 ;
		RECT	8.73 40 8.86 40.05 ;
		RECT	3.02 40.365 3.15 40.415 ;
		RECT	1.57 40.39 1.62 40.52 ;
		RECT	4.87 40.39 4.92 40.52 ;
		RECT	5.9 40.39 5.95 40.52 ;
		RECT	6.375 40.39 6.425 40.52 ;
		RECT	10.27 40.39 10.32 40.52 ;
		RECT	12.65 40.39 12.84 40.52 ;
		RECT	14.33 40.39 14.38 40.52 ;
		RECT	3.02 40.495 3.15 40.545 ;
		RECT	4.035 40.88 4.085 41.01 ;
		RECT	6.835 41.165 6.885 41.215 ;
		RECT	3.02 41.345 3.15 41.395 ;
		RECT	1.57 41.37 1.62 41.5 ;
		RECT	4.87 41.37 4.92 41.5 ;
		RECT	5.9 41.37 5.95 41.5 ;
		RECT	6.375 41.37 6.425 41.5 ;
		RECT	7.015 41.37 7.065 41.5 ;
		RECT	10.27 41.37 10.32 41.5 ;
		RECT	12.79 41.37 12.84 41.5 ;
		RECT	14.33 41.37 14.38 41.5 ;
		RECT	3.02 41.475 3.15 41.525 ;
		RECT	4.035 41.865 4.085 41.995 ;
		RECT	3.02 42.33 3.15 42.38 ;
		RECT	1.57 42.355 1.62 42.485 ;
		RECT	4.87 42.355 4.92 42.485 ;
		RECT	5.9 42.355 5.95 42.485 ;
		RECT	6.375 42.355 6.425 42.485 ;
		RECT	7.015 42.355 7.065 42.485 ;
		RECT	10.27 42.355 10.32 42.485 ;
		RECT	12.79 42.355 12.84 42.485 ;
		RECT	14.33 42.355 14.38 42.485 ;
		RECT	3.02 42.46 3.15 42.51 ;
		RECT	0.9 42.85 0.95 42.98 ;
		RECT	2.485 42.85 2.535 42.98 ;
		RECT	2.615 42.85 2.665 42.98 ;
		RECT	6.065 42.85 6.115 42.98 ;
		RECT	6.675 42.85 6.725 42.98 ;
		RECT	11.555 42.85 11.865 42.98 ;
		RECT	12.52 42.85 12.57 42.98 ;
		RECT	14.005 42.85 14.055 42.98 ;
		RECT	3.8 42.89 3.93 42.94 ;
		RECT	5.635 42.89 5.765 42.94 ;
		RECT	8.31 42.89 8.44 42.94 ;
		RECT	8.73 42.89 8.86 42.94 ;
		RECT	9.315 43.135 9.445 43.185 ;
		RECT	1.045 43.315 1.175 43.365 ;
		RECT	1.34 43.315 1.47 43.365 ;
		RECT	4.47 43.315 4.6 43.365 ;
		RECT	1.86 43.34 1.91 43.47 ;
		RECT	2.01 43.34 2.06 43.47 ;
		RECT	2.32 43.34 2.37 43.47 ;
		RECT	3.25 43.34 3.3 43.47 ;
		RECT	3.515 43.34 3.565 43.47 ;
		RECT	5.035 43.34 5.085 43.47 ;
		RECT	6.22 43.34 6.27 43.47 ;
		RECT	7.5 43.34 7.55 43.47 ;
		RECT	9.72 43.34 9.77 43.47 ;
		RECT	11.025 43.34 11.075 43.47 ;
		RECT	1.045 43.445 1.175 43.495 ;
		RECT	1.34 43.445 1.47 43.495 ;
		RECT	4.47 43.445 4.6 43.495 ;
		RECT	0.62 43.835 0.67 43.965 ;
		RECT	3.65 43.835 3.7 43.965 ;
		RECT	7.19 43.835 7.24 43.965 ;
		RECT	14.14 43.835 14.19 43.965 ;
		RECT	3.02 44.305 3.15 44.355 ;
		RECT	1.57 44.33 1.62 44.46 ;
		RECT	4.87 44.33 4.92 44.46 ;
		RECT	5.9 44.33 5.95 44.46 ;
		RECT	6.375 44.33 6.425 44.46 ;
		RECT	7.015 44.33 7.065 44.46 ;
		RECT	10.27 44.33 10.32 44.46 ;
		RECT	12.79 44.33 12.84 44.46 ;
		RECT	14.335 44.33 14.385 44.46 ;
		RECT	3.02 44.435 3.15 44.485 ;
		RECT	4.035 44.815 4.085 44.945 ;
		RECT	11.685 44.815 11.735 44.945 ;
		RECT	13.9 44.815 13.95 44.945 ;
		RECT	3.02 45.285 3.15 45.335 ;
		RECT	1.57 45.31 1.62 45.44 ;
		RECT	4.87 45.31 4.92 45.44 ;
		RECT	5.9 45.31 5.95 45.44 ;
		RECT	6.375 45.31 6.425 45.44 ;
		RECT	7.015 45.31 7.065 45.44 ;
		RECT	10.27 45.31 10.32 45.44 ;
		RECT	12.79 45.31 12.84 45.44 ;
		RECT	14.335 45.31 14.385 45.44 ;
		RECT	3.02 45.415 3.15 45.465 ;
		RECT	13.8 45.785 13.85 45.915 ;
		RECT	13.675 46.41 13.725 46.54 ;
		RECT	1.085 46.465 1.135 46.595 ;
		RECT	1.38 46.465 1.43 46.595 ;
		RECT	1.86 46.465 1.91 46.595 ;
		RECT	2.01 46.465 2.06 46.595 ;
		RECT	2.32 46.465 2.37 46.595 ;
		RECT	3.25 46.465 3.3 46.595 ;
		RECT	3.515 46.465 3.565 46.595 ;
		RECT	4.51 46.465 4.56 46.595 ;
		RECT	5.035 46.465 5.085 46.595 ;
		RECT	6.22 46.465 6.27 46.595 ;
		RECT	7.5 46.465 7.55 46.595 ;
		RECT	9.72 46.465 9.77 46.595 ;
		RECT	11.025 46.465 11.075 46.595 ;
		RECT	3.8 46.76 3.93 46.81 ;
		RECT	5.635 46.76 5.765 46.81 ;
		RECT	8.31 46.76 8.44 46.81 ;
		RECT	8.73 46.76 8.86 46.81 ;
		RECT	0.9 46.785 0.95 46.915 ;
		RECT	2.485 46.785 2.535 46.915 ;
		RECT	2.615 46.785 2.665 46.915 ;
		RECT	6.065 46.785 6.115 46.915 ;
		RECT	6.675 46.785 6.725 46.915 ;
		RECT	11.555 46.785 11.865 46.915 ;
		RECT	12.52 46.785 12.57 46.915 ;
		RECT	14.005 46.785 14.055 46.915 ;
		RECT	3.8 46.89 3.93 46.94 ;
		RECT	5.635 46.89 5.765 46.94 ;
		RECT	8.31 46.89 8.44 46.94 ;
		RECT	8.73 46.89 8.86 46.94 ;
		RECT	13.9 47.07 13.95 47.12 ;
		RECT	1.045 47.25 1.175 47.3 ;
		RECT	1.34 47.25 1.47 47.3 ;
		RECT	4.47 47.25 4.6 47.3 ;
		RECT	1.86 47.275 1.91 47.405 ;
		RECT	2.01 47.275 2.06 47.405 ;
		RECT	2.32 47.275 2.37 47.405 ;
		RECT	3.25 47.275 3.3 47.405 ;
		RECT	3.515 47.275 3.565 47.405 ;
		RECT	5.035 47.275 5.085 47.405 ;
		RECT	6.22 47.275 6.27 47.405 ;
		RECT	7.5 47.275 7.55 47.405 ;
		RECT	9.72 47.275 9.77 47.405 ;
		RECT	11.025 47.275 11.075 47.405 ;
		RECT	1.045 47.38 1.175 47.43 ;
		RECT	1.34 47.38 1.47 47.43 ;
		RECT	4.47 47.38 4.6 47.43 ;
		RECT	13.9 47.565 13.95 47.615 ;
		RECT	3.8 47.745 3.93 47.795 ;
		RECT	5.635 47.745 5.765 47.795 ;
		RECT	8.31 47.745 8.44 47.795 ;
		RECT	8.73 47.745 8.86 47.795 ;
		RECT	0.9 47.77 0.95 47.9 ;
		RECT	2.485 47.77 2.535 47.9 ;
		RECT	2.615 47.77 2.665 47.9 ;
		RECT	6.065 47.77 6.115 47.9 ;
		RECT	6.675 47.77 6.725 47.9 ;
		RECT	10.12 47.77 10.17 47.9 ;
		RECT	11.555 47.77 11.865 47.9 ;
		RECT	12.52 47.77 12.57 47.9 ;
		RECT	14.005 47.77 14.055 47.9 ;
		RECT	3.8 47.875 3.93 47.925 ;
		RECT	5.635 47.875 5.765 47.925 ;
		RECT	8.31 47.875 8.44 47.925 ;
		RECT	8.73 47.875 8.86 47.925 ;
		RECT	3.02 48.235 3.15 48.285 ;
		RECT	1.57 48.26 1.62 48.39 ;
		RECT	4.87 48.26 4.92 48.39 ;
		RECT	5.9 48.26 5.95 48.39 ;
		RECT	6.375 48.26 6.425 48.39 ;
		RECT	7.015 48.26 7.065 48.39 ;
		RECT	9.11 48.26 9.16 48.39 ;
		RECT	10.27 48.26 10.32 48.39 ;
		RECT	12.79 48.26 12.84 48.39 ;
		RECT	14.335 48.26 14.385 48.39 ;
		RECT	3.02 48.365 3.15 48.415 ;
		RECT	4.035 48.75 4.085 48.88 ;
		RECT	13.9 48.75 13.95 48.88 ;
		RECT	7.19 49.04 7.24 49.09 ;
		RECT	12.655 49.04 12.705 49.09 ;
		RECT	4.035 49.245 4.085 49.375 ;
		RECT	13.9 49.245 13.95 49.375 ;
		RECT	3.02 49.71 3.15 49.76 ;
		RECT	1.57 49.735 1.62 49.865 ;
		RECT	4.87 49.735 4.92 49.865 ;
		RECT	5.9 49.735 5.95 49.865 ;
		RECT	6.375 49.735 6.425 49.865 ;
		RECT	7.015 49.735 7.065 49.865 ;
		RECT	9.11 49.735 9.16 49.865 ;
		RECT	10.27 49.735 10.32 49.865 ;
		RECT	12.79 49.735 12.84 49.865 ;
		RECT	14.335 49.735 14.385 49.865 ;
		RECT	3.02 49.84 3.15 49.89 ;
		RECT	3.8 50.205 3.93 50.255 ;
		RECT	4.22 50.205 4.35 50.255 ;
		RECT	5.635 50.205 5.765 50.255 ;
		RECT	8.31 50.205 8.44 50.255 ;
		RECT	8.73 50.205 8.86 50.255 ;
		RECT	0.9 50.23 0.95 50.36 ;
		RECT	2.485 50.23 2.535 50.36 ;
		RECT	2.615 50.23 2.665 50.36 ;
		RECT	6.065 50.23 6.115 50.36 ;
		RECT	6.675 50.23 6.725 50.36 ;
		RECT	10.12 50.23 10.17 50.36 ;
		RECT	11.555 50.23 11.865 50.36 ;
		RECT	12.52 50.23 12.57 50.36 ;
		RECT	14.005 50.23 14.055 50.36 ;
		RECT	3.8 50.335 3.93 50.385 ;
		RECT	4.22 50.335 4.35 50.385 ;
		RECT	5.635 50.335 5.765 50.385 ;
		RECT	8.31 50.335 8.44 50.385 ;
		RECT	8.73 50.335 8.86 50.385 ;
		RECT	13.9 50.515 13.95 50.565 ;
		RECT	1.045 50.695 1.175 50.745 ;
		RECT	1.34 50.695 1.47 50.745 ;
		RECT	4.47 50.695 4.6 50.745 ;
		RECT	1.86 50.72 1.91 50.85 ;
		RECT	2.01 50.72 2.06 50.85 ;
		RECT	2.32 50.72 2.37 50.85 ;
		RECT	3.25 50.72 3.3 50.85 ;
		RECT	3.515 50.72 3.565 50.85 ;
		RECT	5.035 50.72 5.085 50.85 ;
		RECT	6.22 50.72 6.27 50.85 ;
		RECT	7.5 50.72 7.55 50.85 ;
		RECT	9.72 50.72 9.77 50.85 ;
		RECT	11.025 50.72 11.075 50.85 ;
		RECT	1.045 50.825 1.175 50.875 ;
		RECT	1.34 50.825 1.47 50.875 ;
		RECT	4.47 50.825 4.6 50.875 ;
		RECT	13.9 51.005 13.95 51.055 ;
		RECT	0.9 51.185 14.055 51.365 ;
		RECT	13.675 51.525 13.725 51.655 ;
		RECT	1.085 51.53 1.135 51.66 ;
		RECT	1.38 51.53 1.43 51.66 ;
		RECT	1.86 51.53 1.91 51.66 ;
		RECT	2.01 51.53 2.06 51.66 ;
		RECT	2.32 51.53 2.37 51.66 ;
		RECT	3.25 51.53 3.3 51.66 ;
		RECT	3.515 51.53 3.565 51.66 ;
		RECT	4.51 51.53 4.56 51.66 ;
		RECT	5.035 51.53 5.085 51.66 ;
		RECT	6.22 51.53 6.27 51.66 ;
		RECT	7.5 51.53 7.55 51.66 ;
		RECT	9.72 51.53 9.77 51.66 ;
		RECT	11.025 51.53 11.075 51.66 ;
		RECT	13.8 52.21 13.85 52.34 ;
		RECT	3.02 52.66 3.15 52.71 ;
		RECT	1.57 52.685 1.62 52.815 ;
		RECT	4.87 52.685 4.92 52.815 ;
		RECT	6.375 52.685 6.425 52.815 ;
		RECT	7.015 52.685 7.065 52.815 ;
		RECT	10.27 52.685 10.32 52.815 ;
		RECT	12.79 52.685 12.84 52.815 ;
		RECT	14.33 52.685 14.38 52.815 ;
		RECT	3.02 52.79 3.15 52.84 ;
		RECT	4.035 53.18 4.085 53.31 ;
		RECT	12.655 53.18 12.705 53.31 ;
		RECT	13.9 53.18 13.95 53.31 ;
		RECT	3.02 53.65 3.15 53.7 ;
		RECT	1.57 53.675 1.62 53.805 ;
		RECT	4.87 53.675 4.92 53.805 ;
		RECT	6.375 53.675 6.425 53.805 ;
		RECT	7.015 53.675 7.065 53.805 ;
		RECT	10.27 53.675 10.32 53.805 ;
		RECT	12.79 53.675 12.84 53.805 ;
		RECT	14.33 53.675 14.38 53.805 ;
		RECT	3.02 53.78 3.15 53.83 ;
		RECT	0.62 54.165 0.67 54.295 ;
		RECT	3.65 54.165 3.7 54.295 ;
		RECT	7.19 54.165 7.24 54.295 ;
		RECT	14.14 54.165 14.19 54.295 ;
		RECT	6.85 54.45 6.9 54.5 ;
		RECT	1.045 54.63 1.175 54.68 ;
		RECT	1.34 54.63 1.47 54.68 ;
		RECT	4.47 54.63 4.6 54.68 ;
		RECT	1.86 54.655 1.91 54.785 ;
		RECT	2.01 54.655 2.06 54.785 ;
		RECT	2.32 54.655 2.37 54.785 ;
		RECT	3.25 54.655 3.3 54.785 ;
		RECT	3.515 54.655 3.565 54.785 ;
		RECT	5.035 54.655 5.085 54.785 ;
		RECT	6.22 54.655 6.27 54.785 ;
		RECT	7.5 54.655 7.55 54.785 ;
		RECT	9.72 54.655 9.77 54.785 ;
		RECT	11.025 54.655 11.075 54.785 ;
		RECT	1.045 54.76 1.175 54.81 ;
		RECT	1.34 54.76 1.47 54.81 ;
		RECT	4.47 54.76 4.6 54.81 ;
		RECT	0.9 55.125 14.055 55.305 ;
		RECT	3.02 55.615 3.15 55.665 ;
		RECT	1.57 55.64 1.62 55.77 ;
		RECT	4.87 55.64 4.92 55.77 ;
		RECT	6.375 55.64 6.425 55.77 ;
		RECT	7.015 55.64 7.065 55.77 ;
		RECT	10.27 55.64 10.32 55.77 ;
		RECT	12.79 55.64 12.84 55.77 ;
		RECT	14.33 55.64 14.38 55.77 ;
		RECT	3.02 55.745 3.15 55.795 ;
		RECT	4.035 56.135 4.085 56.265 ;
		RECT	12.655 56.135 12.705 56.265 ;
		RECT	13.9 56.135 13.95 56.265 ;
		RECT	3.02 56.6 3.15 56.65 ;
		RECT	1.57 56.625 1.62 56.755 ;
		RECT	4.87 56.625 4.92 56.755 ;
		RECT	6.375 56.625 6.425 56.755 ;
		RECT	7.015 56.625 7.065 56.755 ;
		RECT	10.27 56.625 10.32 56.755 ;
		RECT	12.79 56.625 12.84 56.755 ;
		RECT	14.33 56.625 14.38 56.755 ;
		RECT	3.02 56.73 3.15 56.78 ;
		RECT	6.85 56.91 6.9 56.96 ;
		RECT	4.035 57.115 4.085 57.245 ;
		RECT	12.655 57.115 12.705 57.245 ;
		RECT	3.02 57.585 3.15 57.635 ;
		RECT	1.57 57.61 1.62 57.74 ;
		RECT	4.87 57.61 4.92 57.74 ;
		RECT	6.375 57.61 6.425 57.74 ;
		RECT	10.27 57.61 10.32 57.74 ;
		RECT	12.79 57.61 12.84 57.74 ;
		RECT	14.33 57.61 14.38 57.74 ;
		RECT	3.02 57.715 3.15 57.765 ;
		RECT	3.8 58.075 3.93 58.125 ;
		RECT	5.635 58.075 5.765 58.125 ;
		RECT	8.31 58.075 8.44 58.125 ;
		RECT	8.73 58.075 8.86 58.125 ;
		RECT	0.9 58.1 0.95 58.23 ;
		RECT	2.485 58.1 2.535 58.23 ;
		RECT	2.615 58.1 2.665 58.23 ;
		RECT	6.065 58.1 6.115 58.23 ;
		RECT	6.725 58.1 6.775 58.23 ;
		RECT	11.555 58.1 12.57 58.23 ;
		RECT	14.005 58.1 14.055 58.23 ;
		RECT	3.8 58.205 3.93 58.255 ;
		RECT	5.635 58.205 5.765 58.255 ;
		RECT	8.31 58.205 8.44 58.255 ;
		RECT	8.73 58.205 8.86 58.255 ;
		RECT	1.045 58.57 1.175 58.62 ;
		RECT	1.34 58.57 1.47 58.62 ;
		RECT	4.47 58.57 4.6 58.62 ;
		RECT	9.275 58.57 9.405 58.62 ;
		RECT	1.86 58.595 1.91 58.725 ;
		RECT	2.01 58.595 2.06 58.725 ;
		RECT	2.32 58.595 2.37 58.725 ;
		RECT	3.25 58.595 3.3 58.725 ;
		RECT	3.515 58.595 3.565 58.725 ;
		RECT	6.22 58.595 6.27 58.725 ;
		RECT	7.5 58.595 7.55 58.725 ;
		RECT	9.72 58.595 9.77 58.725 ;
		RECT	11.025 58.595 11.075 58.725 ;
		RECT	1.045 58.7 1.175 58.75 ;
		RECT	1.34 58.7 1.47 58.75 ;
		RECT	4.47 58.7 4.6 58.75 ;
		RECT	9.275 58.7 9.405 58.75 ;
		RECT	3.8 59.06 3.93 59.11 ;
		RECT	5.635 59.06 5.765 59.11 ;
		RECT	8.31 59.06 8.44 59.11 ;
		RECT	8.73 59.06 8.86 59.11 ;
		RECT	0.9 59.085 0.95 59.215 ;
		RECT	2.485 59.085 2.535 59.215 ;
		RECT	2.615 59.085 2.665 59.215 ;
		RECT	6.065 59.085 6.115 59.215 ;
		RECT	6.725 59.085 6.775 59.215 ;
		RECT	11.555 59.085 11.865 59.215 ;
		RECT	12.52 59.085 12.57 59.215 ;
		RECT	14.005 59.085 14.055 59.215 ;
		RECT	3.8 59.19 3.93 59.24 ;
		RECT	5.635 59.19 5.765 59.24 ;
		RECT	8.31 59.19 8.44 59.24 ;
		RECT	8.73 59.19 8.86 59.24 ;
		RECT	3.02 59.55 3.15 59.6 ;
		RECT	1.57 59.575 1.62 59.705 ;
		RECT	4.87 59.575 4.92 59.705 ;
		RECT	6.375 59.575 6.425 59.705 ;
		RECT	10.27 59.575 10.32 59.705 ;
		RECT	12.79 59.575 12.84 59.705 ;
		RECT	14.33 59.575 14.38 59.705 ;
		RECT	3.02 59.68 3.15 59.73 ;
		RECT	0.9 60.045 14.055 60.225 ;
		RECT	3.02 60.535 3.15 60.585 ;
		RECT	1.57 60.56 1.62 60.69 ;
		RECT	4.87 60.56 4.92 60.69 ;
		RECT	6.375 60.56 6.425 60.69 ;
		RECT	10.27 60.56 10.32 60.69 ;
		RECT	12.79 60.56 12.84 60.69 ;
		RECT	14.33 60.56 14.38 60.69 ;
		RECT	3.02 60.665 3.15 60.715 ;
		RECT	12.655 61.045 12.705 61.175 ;
		RECT	4.035 61.055 4.085 61.185 ;
		RECT	3.02 61.52 3.15 61.57 ;
		RECT	1.57 61.545 1.62 61.675 ;
		RECT	4.87 61.545 4.92 61.675 ;
		RECT	6.375 61.545 6.425 61.675 ;
		RECT	10.27 61.545 10.32 61.675 ;
		RECT	12.79 61.545 12.84 61.675 ;
		RECT	14.33 61.545 14.38 61.675 ;
		RECT	3.02 61.65 3.15 61.7 ;
		RECT	0.9 62.01 14.055 62.19 ;
		RECT	14.29 62.32 14.42 62.37 ;
		RECT	1.045 62.505 1.175 62.555 ;
		RECT	1.34 62.505 1.47 62.555 ;
		RECT	4.47 62.505 4.6 62.555 ;
		RECT	9.275 62.505 9.405 62.555 ;
		RECT	1.86 62.53 1.91 62.66 ;
		RECT	2.01 62.53 2.06 62.66 ;
		RECT	2.32 62.53 2.37 62.66 ;
		RECT	3.25 62.53 3.3 62.66 ;
		RECT	3.515 62.53 3.565 62.66 ;
		RECT	6.22 62.53 6.27 62.66 ;
		RECT	7.5 62.53 7.55 62.66 ;
		RECT	9.72 62.53 9.77 62.66 ;
		RECT	11.025 62.53 11.075 62.66 ;
		RECT	1.045 62.635 1.175 62.685 ;
		RECT	1.34 62.635 1.47 62.685 ;
		RECT	4.47 62.635 4.6 62.685 ;
		RECT	9.275 62.635 9.405 62.685 ;
		RECT	0.9 62.815 0.95 62.865 ;
		RECT	2.51 62.815 2.64 62.865 ;
		RECT	0.9 62.995 14.055 63.175 ;
		RECT	2.18 63.515 2.23 63.645 ;
		RECT	8.56 63.515 8.61 63.645 ;
		RECT	10.27 63.515 10.32 63.645 ;
		RECT	4.035 64.005 4.085 64.135 ;
		RECT	3.02 64.47 3.15 64.52 ;
		RECT	1.57 64.495 1.62 64.625 ;
		RECT	4.87 64.495 4.92 64.625 ;
		RECT	6.375 64.495 6.425 64.625 ;
		RECT	11.69 64.495 11.74 64.625 ;
		RECT	12.79 64.495 12.84 64.625 ;
		RECT	12.79 64.495 12.84 64.625 ;
		RECT	14.33 64.495 14.38 64.625 ;
		RECT	3.02 64.6 3.15 64.65 ;
		RECT	4.035 64.955 4.085 65.085 ;
		RECT	12.655 64.955 12.705 65.085 ;
		RECT	3.02 65.455 3.15 65.505 ;
		RECT	1.57 65.48 1.62 65.61 ;
		RECT	4.87 65.48 4.92 65.61 ;
		RECT	6.375 65.48 6.425 65.61 ;
		RECT	11.69 65.48 11.74 65.61 ;
		RECT	12.79 65.48 12.84 65.61 ;
		RECT	12.79 65.48 12.84 65.61 ;
		RECT	14.33 65.48 14.38 65.61 ;
		RECT	3.02 65.585 3.15 65.635 ;
		RECT	0.9 65.915 14.055 66.095 ;
		RECT	1.045 66.455 1.175 66.505 ;
		RECT	1.34 66.455 1.47 66.505 ;
		RECT	4.47 66.455 4.6 66.505 ;
		RECT	9.275 66.455 9.405 66.505 ;
		RECT	1.86 66.48 1.91 66.61 ;
		RECT	2.01 66.48 2.06 66.61 ;
		RECT	3.25 66.48 3.3 66.61 ;
		RECT	3.515 66.48 3.565 66.61 ;
		RECT	6.22 66.48 6.27 66.61 ;
		RECT	7.5 66.48 7.55 66.61 ;
		RECT	9.72 66.48 9.77 66.61 ;
		RECT	11.025 66.48 11.075 66.61 ;
		RECT	1.045 66.585 1.175 66.635 ;
		RECT	1.34 66.585 1.47 66.635 ;
		RECT	4.47 66.585 4.6 66.635 ;
		RECT	9.275 66.585 9.405 66.635 ;
		RECT	12.655 66.755 12.705 66.805 ;
		RECT	1.045 66.93 1.175 66.98 ;
		RECT	1.34 66.93 1.47 66.98 ;
		RECT	4.47 66.93 4.6 66.98 ;
		RECT	9.275 66.93 9.405 66.98 ;
		RECT	1.86 66.955 1.91 67.085 ;
		RECT	2.01 66.955 2.06 67.085 ;
		RECT	3.25 66.955 3.3 67.085 ;
		RECT	3.515 66.955 3.565 67.085 ;
		RECT	6.22 66.955 6.27 67.085 ;
		RECT	7.5 66.955 7.55 67.085 ;
		RECT	9.72 66.955 9.77 67.085 ;
		RECT	11.025 66.955 11.075 67.085 ;
		RECT	13.675 66.955 13.725 67.085 ;
		RECT	1.045 67.06 1.175 67.11 ;
		RECT	1.34 67.06 1.47 67.11 ;
		RECT	4.47 67.06 4.6 67.11 ;
		RECT	9.275 67.06 9.405 67.11 ;
		RECT	3.02 67.425 3.15 67.475 ;
		RECT	1.57 67.45 1.62 67.58 ;
		RECT	4.87 67.45 4.92 67.58 ;
		RECT	6.375 67.45 6.425 67.58 ;
		RECT	8.975 67.45 9.025 67.58 ;
		RECT	11.69 67.45 11.74 67.58 ;
		RECT	12.79 67.45 12.84 67.58 ;
		RECT	14.33 67.45 14.38 67.58 ;
		RECT	3.02 67.555 3.15 67.605 ;
		RECT	12.655 67.735 12.705 67.785 ;
		RECT	0.9 67.915 14.055 68.095 ;
		RECT	1.57 68.435 1.62 68.565 ;
		RECT	4.87 68.435 4.92 68.565 ;
		RECT	6.375 68.435 6.425 68.565 ;
		RECT	8.975 68.435 9.025 68.565 ;
		RECT	11.69 68.435 11.74 68.565 ;
		RECT	12.79 68.435 12.84 68.565 ;
		RECT	14.33 68.435 14.38 68.565 ;
		RECT	3.02 68.475 3.15 68.525 ;
		RECT	1.045 68.72 1.175 68.77 ;
		RECT	1.34 68.72 1.47 68.77 ;
		RECT	4.47 68.72 4.6 68.77 ;
		RECT	9.275 68.72 9.405 68.77 ;
		RECT	1.86 68.745 1.91 68.875 ;
		RECT	2.01 68.745 2.06 68.875 ;
		RECT	3.25 68.745 3.3 68.875 ;
		RECT	3.515 68.745 3.565 68.875 ;
		RECT	6.22 68.745 6.27 68.875 ;
		RECT	7.5 68.745 7.55 68.875 ;
		RECT	9.72 68.745 9.77 68.875 ;
		RECT	11.025 68.745 11.075 68.875 ;
		RECT	1.045 68.85 1.175 68.9 ;
		RECT	1.34 68.85 1.47 68.9 ;
		RECT	4.47 68.85 4.6 68.9 ;
		RECT	9.275 68.85 9.405 68.9 ;
		RECT	13.8 69.225 13.85 69.355 ;
		RECT	2.18 69.455 2.23 69.585 ;
		RECT	8.56 69.455 8.61 69.585 ;
		RECT	10.27 69.455 10.32 69.585 ;
		RECT	0.62 69.685 0.67 69.815 ;
		RECT	3.65 69.685 3.7 69.815 ;
		RECT	7.19 69.685 7.24 69.815 ;
		RECT	14.14 69.685 14.19 69.815 ;
		RECT	1.085 69.915 1.135 70.045 ;
		RECT	1.38 69.915 1.43 70.045 ;
		RECT	1.86 69.915 1.91 70.045 ;
		RECT	2.01 69.915 2.06 70.045 ;
		RECT	3.25 69.915 3.3 70.045 ;
		RECT	3.515 69.915 3.565 70.045 ;
		RECT	4.51 69.915 4.56 70.045 ;
		RECT	6.22 69.915 6.27 70.045 ;
		RECT	7.5 69.915 7.55 70.045 ;
		RECT	9.315 69.915 9.365 70.045 ;
		RECT	9.72 69.915 9.77 70.045 ;
		RECT	11.025 69.915 11.075 70.045 ;
		RECT	0.435 29.565 0.485 29.695 ;
		RECT	0.435 30.545 0.485 30.675 ;
		RECT	0.435 32.515 0.485 32.645 ;
		RECT	0.435 33.5 0.485 33.63 ;
		RECT	0.435 36.455 0.485 36.585 ;
		RECT	0.435 37.435 0.485 37.565 ;
		RECT	0.435 38.42 0.485 38.55 ;
		RECT	0.435 40.39 0.485 40.52 ;
		RECT	0.17 41.17 0.22 41.22 ;
		RECT	0.435 41.37 0.485 41.5 ;
		RECT	0.435 42.355 0.485 42.485 ;
		RECT	0.18 43.135 0.23 43.185 ;
		RECT	0.435 44.33 0.485 44.46 ;
		RECT	0.435 45.31 0.485 45.44 ;
		RECT	0.435 48.26 0.485 48.39 ;
		RECT	0.435 49.735 0.485 49.865 ;
		RECT	0.435 52.685 0.485 52.815 ;
		RECT	0.435 53.675 0.485 53.805 ;
		RECT	0.18 54.45 0.23 54.5 ;
		RECT	0.435 55.64 0.485 55.77 ;
		RECT	0.435 56.625 0.485 56.755 ;
		RECT	0.17 56.91 0.22 56.96 ;
		RECT	0.435 57.61 0.485 57.74 ;
		RECT	0.435 59.575 0.485 59.705 ;
		RECT	0.435 60.56 0.485 60.69 ;
		RECT	0.435 61.545 0.485 61.675 ;
		RECT	0.17 62.815 0.22 62.865 ;
		RECT	0.435 63.8 0.485 63.85 ;
		RECT	0.435 64.29 0.485 64.34 ;
		RECT	0.435 64.495 0.485 64.625 ;
		RECT	0.435 65.48 0.485 65.61 ;
		RECT	0.435 67.45 0.485 67.58 ;
		RECT	0.435 68.435 0.485 68.565 ;
		RECT	3.06 69.915 3.11 70.045 ;
		RECT	4.87 69.915 4.92 70.045 ;
		RECT	6.375 69.915 6.425 70.045 ;
		RECT	8.975 69.915 9.025 70.045 ;
		RECT	12.79 69.915 12.84 70.045 ;
		RECT	1.57 28.015 1.62 28.145 ;
		RECT	3.06 28.015 3.11 28.145 ;
		RECT	4.87 28.015 4.92 28.145 ;
		RECT	12.79 28.015 12.84 28.145 ;
		RECT	1.57 29.18 1.62 29.31 ;
		RECT	3.02 29.155 3.15 29.335 ;
		RECT	4.87 29.18 4.92 29.31 ;
		RECT	8.955 29.18 9.005 29.31 ;
		RECT	12.79 29.18 12.84 29.31 ;
		RECT	14.29 29.155 14.42 29.335 ;
		RECT	1.045 29.54 1.175 29.72 ;
		RECT	1.34 29.54 1.47 29.72 ;
		RECT	1.86 29.565 1.91 29.695 ;
		RECT	2.01 29.565 2.06 29.695 ;
		RECT	3.25 29.565 3.3 29.695 ;
		RECT	3.515 29.565 3.565 29.695 ;
		RECT	4.47 29.54 4.6 29.72 ;
		RECT	5.035 29.565 5.085 29.695 ;
		RECT	6.22 29.565 6.27 29.695 ;
		RECT	7.5 29.565 7.55 29.695 ;
		RECT	9.275 29.54 9.405 29.72 ;
		RECT	9.72 29.565 9.77 29.695 ;
		RECT	11.025 29.565 11.075 29.695 ;
		RECT	1.045 30.52 1.175 30.7 ;
		RECT	1.34 30.52 1.47 30.7 ;
		RECT	1.86 30.545 1.91 30.675 ;
		RECT	2.01 30.545 2.06 30.675 ;
		RECT	3.25 30.545 3.3 30.675 ;
		RECT	3.515 30.545 3.565 30.675 ;
		RECT	4.47 30.52 4.6 30.7 ;
		RECT	5.035 30.545 5.085 30.675 ;
		RECT	6.22 30.545 6.27 30.675 ;
		RECT	7.5 30.545 7.55 30.675 ;
		RECT	9.275 30.52 9.405 30.7 ;
		RECT	9.72 30.545 9.77 30.675 ;
		RECT	11.025 30.545 11.075 30.675 ;
		RECT	1.57 31.045 1.62 31.175 ;
		RECT	3.02 31.02 3.15 31.2 ;
		RECT	4.87 31.045 4.92 31.175 ;
		RECT	5.9 31.045 5.95 31.175 ;
		RECT	8.955 31.045 9.005 31.175 ;
		RECT	1.57 31.515 1.62 31.645 ;
		RECT	3.02 31.49 3.15 31.67 ;
		RECT	4.87 31.515 4.92 31.645 ;
		RECT	5.9 31.515 5.95 31.645 ;
		RECT	8.955 31.515 9.005 31.645 ;
		RECT	12.79 31.515 12.84 31.645 ;
		RECT	1.045 32.49 1.175 32.67 ;
		RECT	1.34 32.49 1.47 32.67 ;
		RECT	1.86 32.515 1.91 32.645 ;
		RECT	2.01 32.515 2.06 32.645 ;
		RECT	3.25 32.515 3.3 32.645 ;
		RECT	3.515 32.515 3.565 32.645 ;
		RECT	4.47 32.49 4.6 32.67 ;
		RECT	5.035 32.515 5.085 32.645 ;
		RECT	6.22 32.515 6.27 32.645 ;
		RECT	7.5 32.515 7.55 32.645 ;
		RECT	9.275 32.49 9.405 32.67 ;
		RECT	9.72 32.515 9.77 32.645 ;
		RECT	11.025 32.515 11.075 32.645 ;
		RECT	1.045 33.475 1.175 33.655 ;
		RECT	1.34 33.475 1.47 33.655 ;
		RECT	1.86 33.5 1.91 33.63 ;
		RECT	2.01 33.5 2.06 33.63 ;
		RECT	3.25 33.5 3.3 33.63 ;
		RECT	3.515 33.5 3.565 33.63 ;
		RECT	4.47 33.475 4.6 33.655 ;
		RECT	5.035 33.5 5.085 33.63 ;
		RECT	6.22 33.5 6.27 33.63 ;
		RECT	7.5 33.5 7.55 33.63 ;
		RECT	9.72 33.5 9.77 33.63 ;
		RECT	11.025 33.5 11.075 33.63 ;
		RECT	1.57 35.47 1.62 35.6 ;
		RECT	3.02 35.445 3.15 35.625 ;
		RECT	4.87 35.47 4.92 35.6 ;
		RECT	5.9 35.47 5.95 35.6 ;
		RECT	12.79 35.47 12.84 35.6 ;
		RECT	14.29 35.445 14.42 35.625 ;
		RECT	1.045 36.43 1.175 36.61 ;
		RECT	1.34 36.43 1.47 36.61 ;
		RECT	1.86 36.455 1.91 36.585 ;
		RECT	2.01 36.455 2.06 36.585 ;
		RECT	2.32 36.455 2.37 36.585 ;
		RECT	3.25 36.455 3.3 36.585 ;
		RECT	3.515 36.455 3.565 36.585 ;
		RECT	4.47 36.43 4.6 36.61 ;
		RECT	5.035 36.455 5.085 36.585 ;
		RECT	6.22 36.455 6.27 36.585 ;
		RECT	7.5 36.455 7.55 36.585 ;
		RECT	9.72 36.455 9.77 36.585 ;
		RECT	11.025 36.455 11.075 36.585 ;
		RECT	1.045 37.41 1.175 37.59 ;
		RECT	1.34 37.41 1.47 37.59 ;
		RECT	1.86 37.435 1.91 37.565 ;
		RECT	2.01 37.435 2.06 37.565 ;
		RECT	2.32 37.435 2.37 37.565 ;
		RECT	3.25 37.435 3.3 37.565 ;
		RECT	3.515 37.435 3.565 37.565 ;
		RECT	4.47 37.41 4.6 37.59 ;
		RECT	5.035 37.435 5.085 37.565 ;
		RECT	6.22 37.435 6.27 37.565 ;
		RECT	7.5 37.435 7.55 37.565 ;
		RECT	9.72 37.435 9.77 37.565 ;
		RECT	11.025 37.435 11.075 37.565 ;
		RECT	1.045 38.395 1.175 38.575 ;
		RECT	1.34 38.395 1.47 38.575 ;
		RECT	1.86 38.42 1.91 38.55 ;
		RECT	2.01 38.42 2.06 38.55 ;
		RECT	2.32 38.42 2.37 38.55 ;
		RECT	3.25 38.42 3.3 38.55 ;
		RECT	3.515 38.42 3.565 38.55 ;
		RECT	4.47 38.395 4.6 38.575 ;
		RECT	5.035 38.42 5.085 38.55 ;
		RECT	6.22 38.42 6.27 38.55 ;
		RECT	7.5 38.42 7.55 38.55 ;
		RECT	9.72 38.42 9.77 38.55 ;
		RECT	11.025 38.42 11.075 38.55 ;
		RECT	1.57 39.405 1.62 39.535 ;
		RECT	3.02 39.38 3.15 39.56 ;
		RECT	4.87 39.405 4.92 39.535 ;
		RECT	5.9 39.405 5.95 39.535 ;
		RECT	9.43 39.405 9.48 39.535 ;
		RECT	10.27 39.405 10.32 39.535 ;
		RECT	12.79 39.405 12.84 39.535 ;
		RECT	14.29 39.38 14.42 39.56 ;
		RECT	1.045 40.365 1.175 40.545 ;
		RECT	1.34 40.365 1.47 40.545 ;
		RECT	1.86 40.39 1.91 40.52 ;
		RECT	2.01 40.39 2.06 40.52 ;
		RECT	2.32 40.39 2.37 40.52 ;
		RECT	3.25 40.39 3.3 40.52 ;
		RECT	3.515 40.39 3.565 40.52 ;
		RECT	4.47 40.365 4.6 40.545 ;
		RECT	5.035 40.39 5.085 40.52 ;
		RECT	6.22 40.39 6.27 40.52 ;
		RECT	7.5 40.39 7.55 40.52 ;
		RECT	9.72 40.39 9.77 40.52 ;
		RECT	11.025 40.39 11.075 40.52 ;
		RECT	1.045 41.345 1.175 41.525 ;
		RECT	1.34 41.345 1.47 41.525 ;
		RECT	1.86 41.37 1.91 41.5 ;
		RECT	2.01 41.37 2.06 41.5 ;
		RECT	2.32 41.37 2.37 41.5 ;
		RECT	3.25 41.37 3.3 41.5 ;
		RECT	3.515 41.37 3.565 41.5 ;
		RECT	4.47 41.345 4.6 41.525 ;
		RECT	5.035 41.37 5.085 41.5 ;
		RECT	6.22 41.37 6.27 41.5 ;
		RECT	7.5 41.37 7.55 41.5 ;
		RECT	9.72 41.37 9.77 41.5 ;
		RECT	11.025 41.37 11.075 41.5 ;
		RECT	1.045 42.33 1.175 42.51 ;
		RECT	1.34 42.33 1.47 42.51 ;
		RECT	1.86 42.355 1.91 42.485 ;
		RECT	2.01 42.355 2.06 42.485 ;
		RECT	2.32 42.355 2.37 42.485 ;
		RECT	3.25 42.355 3.3 42.485 ;
		RECT	3.515 42.355 3.565 42.485 ;
		RECT	4.47 42.33 4.6 42.51 ;
		RECT	5.035 42.355 5.085 42.485 ;
		RECT	6.22 42.355 6.27 42.485 ;
		RECT	7.5 42.355 7.55 42.485 ;
		RECT	9.72 42.355 9.77 42.485 ;
		RECT	11.025 42.355 11.075 42.485 ;
		RECT	1.57 43.34 1.62 43.47 ;
		RECT	3.02 43.315 3.15 43.495 ;
		RECT	4.87 43.34 4.92 43.47 ;
		RECT	5.9 43.34 5.95 43.47 ;
		RECT	6.375 43.34 6.425 43.47 ;
		RECT	7.015 43.34 7.065 43.47 ;
		RECT	10.27 43.34 10.32 43.47 ;
		RECT	12.79 43.34 12.84 43.47 ;
		RECT	14.29 43.315 14.42 43.495 ;
		RECT	1.045 44.305 1.175 44.485 ;
		RECT	1.34 44.305 1.47 44.485 ;
		RECT	1.86 44.33 1.91 44.46 ;
		RECT	2.01 44.33 2.06 44.46 ;
		RECT	2.32 44.33 2.37 44.46 ;
		RECT	3.25 44.33 3.3 44.46 ;
		RECT	3.515 44.33 3.565 44.46 ;
		RECT	4.47 44.305 4.6 44.485 ;
		RECT	5.035 44.33 5.085 44.46 ;
		RECT	6.22 44.33 6.27 44.46 ;
		RECT	7.5 44.33 7.55 44.46 ;
		RECT	9.72 44.33 9.77 44.46 ;
		RECT	11.025 44.33 11.075 44.46 ;
		RECT	1.045 45.285 1.175 45.465 ;
		RECT	1.34 45.285 1.47 45.465 ;
		RECT	1.86 45.31 1.91 45.44 ;
		RECT	2.01 45.31 2.06 45.44 ;
		RECT	2.32 45.31 2.37 45.44 ;
		RECT	3.25 45.31 3.3 45.44 ;
		RECT	3.515 45.31 3.565 45.44 ;
		RECT	4.47 45.285 4.6 45.465 ;
		RECT	5.035 45.31 5.085 45.44 ;
		RECT	6.22 45.31 6.27 45.44 ;
		RECT	7.5 45.31 7.55 45.44 ;
		RECT	9.72 45.31 9.77 45.44 ;
		RECT	11.025 45.31 11.075 45.44 ;
		RECT	1.57 46.465 1.62 46.595 ;
		RECT	3.06 46.465 3.11 46.595 ;
		RECT	4.87 46.465 4.92 46.595 ;
		RECT	5.9 46.465 5.95 46.595 ;
		RECT	6.375 46.465 6.425 46.595 ;
		RECT	7.015 46.465 7.065 46.595 ;
		RECT	9.11 46.465 9.16 46.595 ;
		RECT	10.27 46.465 10.32 46.595 ;
		RECT	1.57 47.275 1.62 47.405 ;
		RECT	3.02 47.25 3.15 47.43 ;
		RECT	4.87 47.275 4.92 47.405 ;
		RECT	5.9 47.275 5.95 47.405 ;
		RECT	6.375 47.275 6.425 47.405 ;
		RECT	7.015 47.275 7.065 47.405 ;
		RECT	9.11 47.275 9.16 47.405 ;
		RECT	10.27 47.275 10.32 47.405 ;
		RECT	12.79 47.275 12.84 47.405 ;
		RECT	1.045 48.235 1.175 48.415 ;
		RECT	1.34 48.235 1.47 48.415 ;
		RECT	1.86 48.26 1.91 48.39 ;
		RECT	2.01 48.26 2.06 48.39 ;
		RECT	2.32 48.26 2.37 48.39 ;
		RECT	3.25 48.26 3.3 48.39 ;
		RECT	3.515 48.26 3.565 48.39 ;
		RECT	4.47 48.235 4.6 48.415 ;
		RECT	5.035 48.26 5.085 48.39 ;
		RECT	6.22 48.26 6.27 48.39 ;
		RECT	7.5 48.26 7.55 48.39 ;
		RECT	9.72 48.26 9.77 48.39 ;
		RECT	11.025 48.26 11.075 48.39 ;
		RECT	1.045 49.71 1.175 49.89 ;
		RECT	1.34 49.71 1.47 49.89 ;
		RECT	1.86 49.735 1.91 49.865 ;
		RECT	2.01 49.735 2.06 49.865 ;
		RECT	2.32 49.735 2.37 49.865 ;
		RECT	3.25 49.735 3.3 49.865 ;
		RECT	3.515 49.735 3.565 49.865 ;
		RECT	4.47 49.71 4.6 49.89 ;
		RECT	5.035 49.735 5.085 49.865 ;
		RECT	6.22 49.735 6.27 49.865 ;
		RECT	7.5 49.735 7.55 49.865 ;
		RECT	9.72 49.735 9.77 49.865 ;
		RECT	11.025 49.735 11.075 49.865 ;
		RECT	1.57 50.72 1.62 50.85 ;
		RECT	3.02 50.695 3.15 50.875 ;
		RECT	4.87 50.72 4.92 50.85 ;
		RECT	6.375 50.72 6.425 50.85 ;
		RECT	7.015 50.72 7.065 50.85 ;
		RECT	9.11 50.72 9.16 50.85 ;
		RECT	10.27 50.72 10.32 50.85 ;
		RECT	12.79 50.72 12.84 50.85 ;
		RECT	1.57 51.53 1.62 51.66 ;
		RECT	3.06 51.53 3.11 51.66 ;
		RECT	4.87 51.53 4.92 51.66 ;
		RECT	6.375 51.53 6.425 51.66 ;
		RECT	7.015 51.53 7.065 51.66 ;
		RECT	9.11 51.53 9.16 51.66 ;
		RECT	10.27 51.53 10.32 51.66 ;
		RECT	1.045 52.66 1.175 52.84 ;
		RECT	1.34 52.66 1.47 52.84 ;
		RECT	1.86 52.685 1.91 52.815 ;
		RECT	2.01 52.685 2.06 52.815 ;
		RECT	2.32 52.685 2.37 52.815 ;
		RECT	3.25 52.685 3.3 52.815 ;
		RECT	3.515 52.685 3.565 52.815 ;
		RECT	4.47 52.66 4.6 52.84 ;
		RECT	5.035 52.685 5.085 52.815 ;
		RECT	6.22 52.685 6.27 52.815 ;
		RECT	7.5 52.685 7.55 52.815 ;
		RECT	9.72 52.685 9.77 52.815 ;
		RECT	11.025 52.685 11.075 52.815 ;
		RECT	1.045 53.65 1.175 53.83 ;
		RECT	1.34 53.65 1.47 53.83 ;
		RECT	1.86 53.675 1.91 53.805 ;
		RECT	2.01 53.675 2.06 53.805 ;
		RECT	2.32 53.675 2.37 53.805 ;
		RECT	3.25 53.675 3.3 53.805 ;
		RECT	3.515 53.675 3.565 53.805 ;
		RECT	4.47 53.65 4.6 53.83 ;
		RECT	5.035 53.675 5.085 53.805 ;
		RECT	6.22 53.675 6.27 53.805 ;
		RECT	7.5 53.675 7.55 53.805 ;
		RECT	9.72 53.675 9.77 53.805 ;
		RECT	11.025 53.675 11.075 53.805 ;
		RECT	1.57 54.655 1.62 54.785 ;
		RECT	3.02 54.63 3.15 54.81 ;
		RECT	4.87 54.655 4.92 54.785 ;
		RECT	6.375 54.655 6.425 54.785 ;
		RECT	7.015 54.655 7.065 54.785 ;
		RECT	10.27 54.655 10.32 54.785 ;
		RECT	12.79 54.655 12.84 54.785 ;
		RECT	14.29 54.63 14.42 54.81 ;
		RECT	1.045 55.615 1.175 55.795 ;
		RECT	1.34 55.615 1.47 55.795 ;
		RECT	1.86 55.64 1.91 55.77 ;
		RECT	2.01 55.64 2.06 55.77 ;
		RECT	2.32 55.64 2.37 55.77 ;
		RECT	3.25 55.64 3.3 55.77 ;
		RECT	3.515 55.64 3.565 55.77 ;
		RECT	4.47 55.615 4.6 55.795 ;
		RECT	5.035 55.64 5.085 55.77 ;
		RECT	6.22 55.64 6.27 55.77 ;
		RECT	7.5 55.64 7.55 55.77 ;
		RECT	9.275 55.615 9.405 55.795 ;
		RECT	9.72 55.64 9.77 55.77 ;
		RECT	11.025 55.64 11.075 55.77 ;
		RECT	1.045 56.6 1.175 56.78 ;
		RECT	1.34 56.6 1.47 56.78 ;
		RECT	1.86 56.625 1.91 56.755 ;
		RECT	2.01 56.625 2.06 56.755 ;
		RECT	2.32 56.625 2.37 56.755 ;
		RECT	3.25 56.625 3.3 56.755 ;
		RECT	3.515 56.625 3.565 56.755 ;
		RECT	4.47 56.6 4.6 56.78 ;
		RECT	5.035 56.625 5.085 56.755 ;
		RECT	6.22 56.625 6.27 56.755 ;
		RECT	7.5 56.625 7.55 56.755 ;
		RECT	9.275 56.6 9.405 56.78 ;
		RECT	9.72 56.625 9.77 56.755 ;
		RECT	11.025 56.625 11.075 56.755 ;
		RECT	1.045 57.585 1.175 57.765 ;
		RECT	1.34 57.585 1.47 57.765 ;
		RECT	1.86 57.61 1.91 57.74 ;
		RECT	2.01 57.61 2.06 57.74 ;
		RECT	2.32 57.61 2.37 57.74 ;
		RECT	3.25 57.61 3.3 57.74 ;
		RECT	3.515 57.61 3.565 57.74 ;
		RECT	4.47 57.585 4.6 57.765 ;
		RECT	6.22 57.61 6.27 57.74 ;
		RECT	7.5 57.61 7.55 57.74 ;
		RECT	9.275 57.585 9.405 57.765 ;
		RECT	9.72 57.61 9.77 57.74 ;
		RECT	11.025 57.61 11.075 57.74 ;
		RECT	1.57 58.595 1.62 58.725 ;
		RECT	3.02 58.57 3.15 58.75 ;
		RECT	4.87 58.595 4.92 58.725 ;
		RECT	6.375 58.595 6.425 58.725 ;
		RECT	10 58.595 10.05 58.725 ;
		RECT	10.27 58.595 10.32 58.725 ;
		RECT	12.79 58.595 12.84 58.725 ;
		RECT	14.29 58.57 14.42 58.75 ;
		RECT	1.045 59.55 1.175 59.73 ;
		RECT	1.34 59.55 1.47 59.73 ;
		RECT	1.86 59.575 1.91 59.705 ;
		RECT	2.01 59.575 2.06 59.705 ;
		RECT	2.32 59.575 2.37 59.705 ;
		RECT	3.25 59.575 3.3 59.705 ;
		RECT	3.515 59.575 3.565 59.705 ;
		RECT	4.47 59.55 4.6 59.73 ;
		RECT	6.22 59.575 6.27 59.705 ;
		RECT	7.5 59.575 7.55 59.705 ;
		RECT	9.275 59.55 9.405 59.73 ;
		RECT	9.72 59.575 9.77 59.705 ;
		RECT	11.025 59.575 11.075 59.705 ;
		RECT	1.045 60.535 1.175 60.715 ;
		RECT	1.34 60.535 1.47 60.715 ;
		RECT	1.86 60.56 1.91 60.69 ;
		RECT	2.01 60.56 2.06 60.69 ;
		RECT	2.32 60.56 2.37 60.69 ;
		RECT	3.25 60.56 3.3 60.69 ;
		RECT	3.515 60.56 3.565 60.69 ;
		RECT	4.47 60.535 4.6 60.715 ;
		RECT	6.22 60.56 6.27 60.69 ;
		RECT	7.5 60.56 7.55 60.69 ;
		RECT	9.275 60.535 9.405 60.715 ;
		RECT	9.72 60.56 9.77 60.69 ;
		RECT	11.025 60.56 11.075 60.69 ;
		RECT	1.045 61.52 1.175 61.7 ;
		RECT	1.34 61.52 1.47 61.7 ;
		RECT	1.86 61.545 1.91 61.675 ;
		RECT	2.01 61.545 2.06 61.675 ;
		RECT	2.32 61.545 2.37 61.675 ;
		RECT	3.25 61.545 3.3 61.675 ;
		RECT	3.515 61.545 3.565 61.675 ;
		RECT	4.47 61.52 4.6 61.7 ;
		RECT	6.22 61.545 6.27 61.675 ;
		RECT	7.5 61.545 7.55 61.675 ;
		RECT	9.275 61.52 9.405 61.7 ;
		RECT	9.72 61.545 9.77 61.675 ;
		RECT	11.025 61.545 11.075 61.675 ;
		RECT	1.57 62.53 1.62 62.66 ;
		RECT	3.02 62.505 3.15 62.685 ;
		RECT	4.87 62.53 4.92 62.66 ;
		RECT	6.375 62.53 6.425 62.66 ;
		RECT	12.79 62.53 12.84 62.66 ;
		RECT	14.29 62.505 14.42 62.685 ;
		RECT	1.045 64.47 1.175 64.65 ;
		RECT	1.34 64.47 1.47 64.65 ;
		RECT	1.86 64.495 1.91 64.625 ;
		RECT	2.01 64.495 2.06 64.625 ;
		RECT	2.32 64.495 2.37 64.625 ;
		RECT	3.25 64.495 3.3 64.625 ;
		RECT	3.515 64.495 3.565 64.625 ;
		RECT	4.47 64.47 4.6 64.65 ;
		RECT	6.22 64.495 6.27 64.625 ;
		RECT	7.5 64.495 7.55 64.625 ;
		RECT	9.275 64.47 9.405 64.65 ;
		RECT	9.72 64.495 9.77 64.625 ;
		RECT	11.025 64.495 11.075 64.625 ;
		RECT	1.045 65.455 1.175 65.635 ;
		RECT	1.34 65.455 1.47 65.635 ;
		RECT	1.86 65.48 1.91 65.61 ;
		RECT	2.01 65.48 2.06 65.61 ;
		RECT	2.32 65.48 2.37 65.61 ;
		RECT	3.25 65.48 3.3 65.61 ;
		RECT	3.515 65.48 3.565 65.61 ;
		RECT	4.47 65.455 4.6 65.635 ;
		RECT	6.22 65.48 6.27 65.61 ;
		RECT	7.5 65.48 7.55 65.61 ;
		RECT	9.275 65.455 9.405 65.635 ;
		RECT	9.72 65.48 9.77 65.61 ;
		RECT	11.025 65.48 11.075 65.61 ;
		RECT	1.57 66.48 1.62 66.61 ;
		RECT	3.02 66.455 3.15 66.635 ;
		RECT	4.87 66.48 4.92 66.61 ;
		RECT	6.375 66.48 6.425 66.61 ;
		RECT	11.69 66.48 11.74 66.61 ;
		RECT	12.79 66.48 12.84 66.61 ;
		RECT	1.57 66.955 1.62 67.085 ;
		RECT	3.02 66.93 3.15 67.11 ;
		RECT	4.87 66.955 4.92 67.085 ;
		RECT	6.375 66.955 6.425 67.085 ;
		RECT	1.045 67.425 1.175 67.605 ;
		RECT	1.34 67.425 1.47 67.605 ;
		RECT	1.86 67.45 1.91 67.58 ;
		RECT	2.01 67.45 2.06 67.58 ;
		RECT	3.25 67.45 3.3 67.58 ;
		RECT	3.515 67.45 3.565 67.58 ;
		RECT	4.47 67.425 4.6 67.605 ;
		RECT	6.22 67.45 6.27 67.58 ;
		RECT	7.5 67.45 7.55 67.58 ;
		RECT	9.275 67.425 9.405 67.605 ;
		RECT	9.72 67.45 9.77 67.58 ;
		RECT	11.025 67.45 11.075 67.58 ;
		RECT	1.86 68.435 1.91 68.565 ;
		RECT	2.01 68.435 2.06 68.565 ;
		RECT	3.25 68.435 3.3 68.565 ;
		RECT	3.515 68.435 3.565 68.565 ;
		RECT	6.22 68.435 6.27 68.565 ;
		RECT	7.5 68.435 7.55 68.565 ;
		RECT	9.72 68.435 9.77 68.565 ;
		RECT	11.025 68.435 11.075 68.565 ;
		RECT	1.57 68.745 1.62 68.875 ;
		RECT	3.02 68.72 3.15 68.9 ;
		RECT	4.87 68.745 4.92 68.875 ;
		RECT	6.375 68.745 6.425 68.875 ;
		RECT	8.975 68.745 9.025 68.875 ;
		RECT	12.79 68.745 12.84 68.875 ;
		RECT	14.29 68.72 14.42 68.9 ;
		RECT	0.9 28.245 0.95 28.375 ;
		RECT	2.485 28.245 2.665 28.375 ;
		RECT	3.84 28.245 3.89 28.375 ;
		RECT	5.675 28.245 5.725 28.375 ;
		RECT	6.065 28.245 6.115 28.375 ;
		RECT	6.725 28.245 6.775 28.375 ;
		RECT	8.35 28.245 8.4 28.375 ;
		RECT	8.77 28.245 8.82 28.375 ;
		RECT	11.555 28.245 11.605 28.375 ;
		RECT	11.815 28.245 11.865 28.375 ;
		RECT	12.52 28.245 12.57 28.375 ;
		RECT	14.005 28.245 14.055 28.375 ;
		RECT	0.62 30.055 0.67 30.185 ;
		RECT	3.65 30.055 3.7 30.185 ;
		RECT	7.18 30.055 7.23 30.185 ;
		RECT	14.14 30.055 14.19 30.185 ;
		RECT	0.62 32.06 0.67 32.19 ;
		RECT	3.65 32.06 3.7 32.19 ;
		RECT	7.18 32.06 7.23 32.19 ;
		RECT	14.14 32.06 14.19 32.19 ;
		RECT	0.62 34.975 0.67 35.105 ;
		RECT	3.65 34.975 3.7 35.105 ;
		RECT	7.18 34.975 7.23 35.105 ;
		RECT	14.14 34.975 14.19 35.105 ;
		RECT	0.62 35.96 0.67 36.09 ;
		RECT	3.65 35.96 3.7 36.09 ;
		RECT	7.18 35.96 7.23 36.09 ;
		RECT	14.14 35.96 14.19 36.09 ;
		RECT	0.62 37.93 0.67 38.06 ;
		RECT	3.65 37.93 3.7 38.06 ;
		RECT	7.18 37.93 7.23 38.06 ;
		RECT	14.14 37.93 14.19 38.06 ;
		RECT	0.62 38.91 0.67 39.04 ;
		RECT	3.65 38.91 3.7 39.04 ;
		RECT	7.18 38.91 7.23 39.04 ;
		RECT	14.14 38.91 14.19 39.04 ;
		RECT	0.62 39.895 0.67 40.025 ;
		RECT	3.65 39.895 3.7 40.025 ;
		RECT	7.18 39.895 7.23 40.025 ;
		RECT	14.14 39.895 14.19 40.025 ;
		RECT	0.62 42.85 0.67 42.98 ;
		RECT	3.65 42.85 3.7 42.98 ;
		RECT	7.18 42.85 7.23 42.98 ;
		RECT	14.14 42.85 14.19 42.98 ;
		RECT	0.9 43.835 0.95 43.965 ;
		RECT	2.485 43.835 2.665 43.965 ;
		RECT	3.8 43.81 3.93 43.99 ;
		RECT	5.635 43.81 5.765 43.99 ;
		RECT	6.065 43.835 6.115 43.965 ;
		RECT	6.675 43.835 6.725 43.965 ;
		RECT	8.31 43.81 8.44 43.99 ;
		RECT	8.73 43.81 8.86 43.99 ;
		RECT	11.555 43.835 11.605 43.965 ;
		RECT	11.815 43.835 11.865 43.965 ;
		RECT	12.52 43.835 12.57 43.965 ;
		RECT	14.005 43.835 14.055 43.965 ;
		RECT	0.62 46.785 0.67 46.915 ;
		RECT	3.65 46.785 3.7 46.915 ;
		RECT	7.18 46.785 7.23 46.915 ;
		RECT	14.14 46.785 14.19 46.915 ;
		RECT	0.62 47.77 0.67 47.9 ;
		RECT	3.65 47.77 3.7 47.9 ;
		RECT	7.18 47.77 7.23 47.9 ;
		RECT	14.14 47.77 14.19 47.9 ;
		RECT	8.31 49.04 8.44 49.09 ;
		RECT	8.73 49.04 8.86 49.09 ;
		RECT	10.12 49.04 10.17 49.09 ;
		RECT	11.555 49.04 11.605 49.09 ;
		RECT	11.815 49.04 11.865 49.09 ;
		RECT	12.52 49.04 12.57 49.09 ;
		RECT	0.62 50.23 0.67 50.36 ;
		RECT	3.65 50.23 3.7 50.36 ;
		RECT	7.18 50.23 7.23 50.36 ;
		RECT	12.655 50.23 12.705 50.36 ;
		RECT	14.14 50.23 14.19 50.36 ;
		RECT	0.62 51.21 0.67 51.34 ;
		RECT	3.65 51.21 3.7 51.34 ;
		RECT	7.18 51.21 7.23 51.34 ;
		RECT	14.14 51.21 14.19 51.34 ;
		RECT	0.9 54.165 0.95 54.295 ;
		RECT	2.51 54.14 2.64 54.32 ;
		RECT	3.8 54.14 3.93 54.32 ;
		RECT	5.635 54.14 5.765 54.32 ;
		RECT	6.065 54.165 6.115 54.295 ;
		RECT	6.675 54.165 6.725 54.295 ;
		RECT	8.31 54.14 8.44 54.32 ;
		RECT	8.73 54.14 8.86 54.32 ;
		RECT	11.555 54.165 11.605 54.295 ;
		RECT	11.815 54.165 11.865 54.295 ;
		RECT	12.52 54.165 12.57 54.295 ;
		RECT	14.005 54.165 14.055 54.295 ;
		RECT	0.62 55.15 0.67 55.28 ;
		RECT	3.65 55.15 3.7 55.28 ;
		RECT	7.18 55.15 7.23 55.28 ;
		RECT	14.14 55.15 14.19 55.28 ;
		RECT	0.62 58.1 0.67 58.23 ;
		RECT	3.65 58.1 3.7 58.23 ;
		RECT	7.18 58.1 7.23 58.23 ;
		RECT	14.14 58.1 14.19 58.23 ;
		RECT	0.62 59.085 0.67 59.215 ;
		RECT	3.65 59.085 3.7 59.215 ;
		RECT	7.18 59.085 7.23 59.215 ;
		RECT	14.14 59.085 14.19 59.215 ;
		RECT	0.62 60.07 0.67 60.2 ;
		RECT	3.65 60.07 3.7 60.2 ;
		RECT	7.18 60.07 7.23 60.2 ;
		RECT	14.14 60.07 14.19 60.2 ;
		RECT	0.62 62.035 0.67 62.165 ;
		RECT	3.65 62.035 3.7 62.165 ;
		RECT	7.18 62.035 7.23 62.165 ;
		RECT	14.14 62.035 14.19 62.165 ;
		RECT	0.62 62.815 0.67 62.865 ;
		RECT	0.62 63.02 0.67 63.15 ;
		RECT	3.65 63.02 3.7 63.15 ;
		RECT	7.18 63.02 7.23 63.15 ;
		RECT	14.14 63.02 14.19 63.15 ;
		RECT	0.62 65.94 0.67 66.07 ;
		RECT	3.65 65.94 3.7 66.07 ;
		RECT	7.18 65.94 7.23 66.07 ;
		RECT	14.14 65.94 14.19 66.07 ;
		RECT	0.62 67.94 0.67 68.07 ;
		RECT	3.65 67.94 3.7 68.07 ;
		RECT	7.18 67.94 7.23 68.07 ;
		RECT	14.14 67.94 14.19 68.07 ;
		RECT	0.9 69.685 0.95 69.815 ;
		RECT	2.485 69.685 2.665 69.815 ;
		RECT	3.84 69.685 3.89 69.815 ;
		RECT	5.675 69.685 5.725 69.815 ;
		RECT	6.065 69.685 6.115 69.815 ;
		RECT	6.725 69.685 6.775 69.815 ;
		RECT	8.35 69.685 8.4 69.815 ;
		RECT	8.77 69.685 8.82 69.815 ;
		RECT	11.555 69.685 11.605 69.815 ;
		RECT	11.815 69.685 11.865 69.815 ;
		RECT	12.52 69.685 12.57 69.815 ;
		RECT	14.005 69.685 14.055 69.815 ;
		RECT	1.57 28.475 1.62 28.605 ;
		RECT	3.06 28.475 3.11 28.605 ;
		RECT	4.87 28.475 4.92 28.605 ;
		RECT	12.79 28.475 12.84 28.605 ;
		RECT	14.33 28.475 14.38 28.605 ;
		RECT	2.18 29.565 2.23 29.695 ;
		RECT	8.56 29.565 8.61 29.695 ;
		RECT	10.27 29.565 10.32 29.695 ;
		RECT	2.18 30.545 2.23 30.675 ;
		RECT	8.56 30.545 8.61 30.675 ;
		RECT	10.27 30.545 10.32 30.675 ;
		RECT	2.18 32.515 2.23 32.645 ;
		RECT	8.56 32.515 8.61 32.645 ;
		RECT	10.27 32.515 10.32 32.645 ;
		RECT	2.18 33.5 2.23 33.63 ;
		RECT	8.56 33.5 8.61 33.63 ;
		RECT	10.27 33.5 10.32 33.63 ;
		RECT	1.57 34.485 1.62 34.615 ;
		RECT	3.02 34.46 3.15 34.64 ;
		RECT	4.87 34.485 4.92 34.615 ;
		RECT	5.9 34.485 5.95 34.615 ;
		RECT	12.79 34.485 12.84 34.615 ;
		RECT	14.29 34.46 14.42 34.64 ;
		RECT	2.18 36.455 2.23 36.585 ;
		RECT	8.56 36.455 8.61 36.585 ;
		RECT	2.18 37.435 2.23 37.565 ;
		RECT	8.56 37.435 8.61 37.565 ;
		RECT	2.18 38.42 2.23 38.55 ;
		RECT	8.56 38.42 8.61 38.55 ;
		RECT	2.18 40.39 2.23 40.52 ;
		RECT	8.56 40.39 8.61 40.52 ;
		RECT	2.18 41.37 2.23 41.5 ;
		RECT	8.56 41.37 8.61 41.5 ;
		RECT	2.18 42.355 2.23 42.485 ;
		RECT	8.56 42.355 8.61 42.485 ;
		RECT	2.18 44.33 2.23 44.46 ;
		RECT	8.56 44.33 8.61 44.46 ;
		RECT	2.18 45.31 2.23 45.44 ;
		RECT	8.56 45.31 8.61 45.44 ;
		RECT	2.18 48.26 2.23 48.39 ;
		RECT	8.56 48.26 8.61 48.39 ;
		RECT	2.18 49.735 2.23 49.865 ;
		RECT	8.56 49.735 8.61 49.865 ;
		RECT	2.18 52.685 2.23 52.815 ;
		RECT	8.56 52.685 8.61 52.815 ;
		RECT	2.18 53.675 2.23 53.805 ;
		RECT	8.56 53.675 8.61 53.805 ;
		RECT	2.18 55.64 2.23 55.77 ;
		RECT	8.56 55.64 8.61 55.77 ;
		RECT	2.18 56.625 2.23 56.755 ;
		RECT	8.56 56.625 8.61 56.755 ;
		RECT	2.18 57.61 2.23 57.74 ;
		RECT	8.56 57.61 8.61 57.74 ;
		RECT	2.18 59.575 2.23 59.705 ;
		RECT	8.56 59.575 8.61 59.705 ;
		RECT	2.18 60.56 2.23 60.69 ;
		RECT	8.56 60.56 8.61 60.69 ;
		RECT	2.18 61.545 2.23 61.675 ;
		RECT	8.56 61.545 8.61 61.675 ;
		RECT	1.57 63.515 1.62 63.645 ;
		RECT	3.02 63.49 3.15 63.67 ;
		RECT	4.87 63.515 4.92 63.645 ;
		RECT	6.375 63.515 6.425 63.645 ;
		RECT	12.79 63.515 12.84 63.645 ;
		RECT	14.29 63.49 14.42 63.67 ;
		RECT	2.18 64.495 2.23 64.625 ;
		RECT	8.56 64.495 8.61 64.625 ;
		RECT	10.27 64.495 10.32 64.625 ;
		RECT	2.18 65.48 2.23 65.61 ;
		RECT	8.56 65.48 8.61 65.61 ;
		RECT	10.27 65.48 10.32 65.61 ;
		RECT	2.18 67.45 2.23 67.58 ;
		RECT	8.56 67.45 8.61 67.58 ;
		RECT	10.27 67.45 10.32 67.58 ;
		RECT	2.18 68.435 2.23 68.565 ;
		RECT	8.56 68.435 8.61 68.565 ;
		RECT	10.27 68.435 10.32 68.565 ;
		RECT	3.06 69.455 3.11 69.585 ;
		RECT	4.87 69.455 4.92 69.585 ;
		RECT	6.375 69.455 6.425 69.585 ;
		RECT	8.975 69.455 9.025 69.585 ;
		RECT	12.79 69.455 12.84 69.585 ;
		RECT	14.33 69.455 14.38 69.585 ;
		RECT	20.875 0.425 21.055 0.555 ;
		RECT	14.965 0.655 15.015 0.785 ;
		RECT	19.485 0.655 19.535 0.785 ;
		RECT	14.765 0.655 14.815 0.785 ;
		RECT	19.685 0.655 19.735 0.785 ;
		RECT	20.7 0.425 20.75 0.555 ;
		RECT	20.875 100.385 21.055 100.515 ;
		RECT	14.965 100.155 15.015 100.285 ;
		RECT	19.485 100.155 19.535 100.285 ;
		RECT	14.765 100.155 14.815 100.285 ;
		RECT	19.685 100.155 19.735 100.285 ;
		RECT	20.7 100.385 20.75 100.515 ;
		RECT	14.565 3.305 14.615 3.435 ;
		RECT	19.885 3.305 19.935 3.435 ;
		RECT	14.765 3.535 14.815 3.665 ;
		RECT	14.765 1.115 14.815 1.245 ;
		RECT	19.685 3.535 19.735 3.665 ;
		RECT	19.685 1.115 19.735 1.245 ;
		RECT	14.965 3.535 15.015 3.665 ;
		RECT	14.965 1.115 15.015 1.245 ;
		RECT	19.485 3.535 19.535 3.665 ;
		RECT	19.485 1.115 19.535 1.245 ;
		RECT	14.565 26.345 14.615 26.475 ;
		RECT	19.885 26.345 19.935 26.475 ;
		RECT	14.765 26.575 14.815 26.705 ;
		RECT	14.765 24.155 14.815 24.285 ;
		RECT	19.685 26.575 19.735 26.705 ;
		RECT	19.685 24.155 19.735 24.285 ;
		RECT	14.965 26.575 15.015 26.705 ;
		RECT	14.965 24.155 15.015 24.285 ;
		RECT	19.485 26.575 19.535 26.705 ;
		RECT	19.485 24.155 19.535 24.285 ;
		RECT	14.565 23.465 14.615 23.595 ;
		RECT	19.885 23.465 19.935 23.595 ;
		RECT	14.765 23.695 14.815 23.825 ;
		RECT	14.765 21.275 14.815 21.405 ;
		RECT	19.685 23.695 19.735 23.825 ;
		RECT	19.685 21.275 19.735 21.405 ;
		RECT	14.965 23.695 15.015 23.825 ;
		RECT	14.965 21.275 15.015 21.405 ;
		RECT	19.485 23.695 19.535 23.825 ;
		RECT	19.485 21.275 19.535 21.405 ;
		RECT	14.565 20.585 14.615 20.715 ;
		RECT	19.885 20.585 19.935 20.715 ;
		RECT	14.765 20.815 14.815 20.945 ;
		RECT	14.765 18.395 14.815 18.525 ;
		RECT	19.685 20.815 19.735 20.945 ;
		RECT	19.685 18.395 19.735 18.525 ;
		RECT	14.965 20.815 15.015 20.945 ;
		RECT	14.965 18.395 15.015 18.525 ;
		RECT	19.485 20.815 19.535 20.945 ;
		RECT	19.485 18.395 19.535 18.525 ;
		RECT	14.565 17.705 14.615 17.835 ;
		RECT	19.885 17.705 19.935 17.835 ;
		RECT	14.765 17.935 14.815 18.065 ;
		RECT	14.765 15.515 14.815 15.645 ;
		RECT	19.685 17.935 19.735 18.065 ;
		RECT	19.685 15.515 19.735 15.645 ;
		RECT	14.965 17.935 15.015 18.065 ;
		RECT	14.965 15.515 15.015 15.645 ;
		RECT	19.485 17.935 19.535 18.065 ;
		RECT	19.485 15.515 19.535 15.645 ;
		RECT	14.565 14.825 14.615 14.955 ;
		RECT	19.885 14.825 19.935 14.955 ;
		RECT	14.765 15.055 14.815 15.185 ;
		RECT	14.765 12.635 14.815 12.765 ;
		RECT	19.685 15.055 19.735 15.185 ;
		RECT	19.685 12.635 19.735 12.765 ;
		RECT	14.965 15.055 15.015 15.185 ;
		RECT	14.965 12.635 15.015 12.765 ;
		RECT	19.485 15.055 19.535 15.185 ;
		RECT	19.485 12.635 19.535 12.765 ;
		RECT	14.565 11.945 14.615 12.075 ;
		RECT	19.885 11.945 19.935 12.075 ;
		RECT	14.765 12.175 14.815 12.305 ;
		RECT	14.765 9.755 14.815 9.885 ;
		RECT	19.685 12.175 19.735 12.305 ;
		RECT	19.685 9.755 19.735 9.885 ;
		RECT	14.965 12.175 15.015 12.305 ;
		RECT	14.965 9.755 15.015 9.885 ;
		RECT	19.485 12.175 19.535 12.305 ;
		RECT	19.485 9.755 19.535 9.885 ;
		RECT	14.565 9.065 14.615 9.195 ;
		RECT	19.885 9.065 19.935 9.195 ;
		RECT	14.765 9.295 14.815 9.425 ;
		RECT	14.765 6.875 14.815 7.005 ;
		RECT	19.685 9.295 19.735 9.425 ;
		RECT	19.685 6.875 19.735 7.005 ;
		RECT	14.965 9.295 15.015 9.425 ;
		RECT	14.965 6.875 15.015 7.005 ;
		RECT	19.485 9.295 19.535 9.425 ;
		RECT	19.485 6.875 19.535 7.005 ;
		RECT	14.565 6.185 14.615 6.315 ;
		RECT	19.885 6.185 19.935 6.315 ;
		RECT	14.765 6.415 14.815 6.545 ;
		RECT	14.765 3.995 14.815 4.125 ;
		RECT	19.685 6.415 19.735 6.545 ;
		RECT	19.685 3.995 19.735 4.125 ;
		RECT	14.965 6.415 15.015 6.545 ;
		RECT	14.965 3.995 15.015 4.125 ;
		RECT	19.485 6.415 19.535 6.545 ;
		RECT	19.485 3.995 19.535 4.125 ;
		RECT	20.085 23.695 20.265 23.825 ;
		RECT	20.875 23.465 21.055 23.595 ;
		RECT	20.085 21.275 20.265 21.405 ;
		RECT	20.43 21.045 20.48 21.175 ;
		RECT	20.085 20.815 20.265 20.945 ;
		RECT	20.875 20.585 21.055 20.715 ;
		RECT	20.085 18.395 20.265 18.525 ;
		RECT	20.43 18.165 20.48 18.295 ;
		RECT	20.085 17.935 20.265 18.065 ;
		RECT	20.875 17.705 21.055 17.835 ;
		RECT	20.085 15.515 20.265 15.645 ;
		RECT	20.43 15.285 20.48 15.415 ;
		RECT	20.085 15.055 20.265 15.185 ;
		RECT	20.875 14.825 21.055 14.955 ;
		RECT	20.085 12.635 20.265 12.765 ;
		RECT	20.43 12.405 20.48 12.535 ;
		RECT	20.085 12.175 20.265 12.305 ;
		RECT	20.875 11.945 21.055 12.075 ;
		RECT	20.085 9.755 20.265 9.885 ;
		RECT	20.43 9.525 20.48 9.655 ;
		RECT	20.085 9.295 20.265 9.425 ;
		RECT	20.875 9.065 21.055 9.195 ;
		RECT	20.085 6.875 20.265 7.005 ;
		RECT	20.43 6.645 20.48 6.775 ;
		RECT	20.085 6.415 20.265 6.545 ;
		RECT	20.875 6.185 21.055 6.315 ;
		RECT	20.085 3.995 20.265 4.125 ;
		RECT	20.43 3.765 20.48 3.895 ;
		RECT	20.085 3.535 20.265 3.665 ;
		RECT	20.875 3.305 21.055 3.435 ;
		RECT	20.085 1.115 20.265 1.245 ;
		RECT	20.43 0.885 20.48 1.015 ;
		RECT	20.085 26.575 20.265 26.705 ;
		RECT	20.875 26.345 21.055 26.475 ;
		RECT	20.085 24.155 20.265 24.285 ;
		RECT	20.43 23.925 20.48 24.055 ;
		RECT	14.565 97.505 14.615 97.635 ;
		RECT	19.885 97.505 19.935 97.635 ;
		RECT	14.765 97.275 14.815 97.405 ;
		RECT	14.765 99.695 14.815 99.825 ;
		RECT	19.685 97.275 19.735 97.405 ;
		RECT	19.685 99.695 19.735 99.825 ;
		RECT	14.965 97.275 15.015 97.405 ;
		RECT	14.965 99.695 15.015 99.825 ;
		RECT	19.485 97.275 19.535 97.405 ;
		RECT	19.485 99.695 19.535 99.825 ;
		RECT	14.565 71.585 14.615 71.715 ;
		RECT	19.885 71.585 19.935 71.715 ;
		RECT	14.765 71.355 14.815 71.485 ;
		RECT	14.765 73.775 14.815 73.905 ;
		RECT	19.685 71.355 19.735 71.485 ;
		RECT	19.685 73.775 19.735 73.905 ;
		RECT	14.965 71.355 15.015 71.485 ;
		RECT	14.965 73.775 15.015 73.905 ;
		RECT	19.485 71.355 19.535 71.485 ;
		RECT	19.485 73.775 19.535 73.905 ;
		RECT	14.565 74.465 14.615 74.595 ;
		RECT	19.885 74.465 19.935 74.595 ;
		RECT	14.765 74.235 14.815 74.365 ;
		RECT	14.765 76.655 14.815 76.785 ;
		RECT	19.685 74.235 19.735 74.365 ;
		RECT	19.685 76.655 19.735 76.785 ;
		RECT	14.965 74.235 15.015 74.365 ;
		RECT	14.965 76.655 15.015 76.785 ;
		RECT	19.485 74.235 19.535 74.365 ;
		RECT	19.485 76.655 19.535 76.785 ;
		RECT	14.565 77.345 14.615 77.475 ;
		RECT	19.885 77.345 19.935 77.475 ;
		RECT	14.765 77.115 14.815 77.245 ;
		RECT	14.765 79.535 14.815 79.665 ;
		RECT	19.685 77.115 19.735 77.245 ;
		RECT	19.685 79.535 19.735 79.665 ;
		RECT	14.965 77.115 15.015 77.245 ;
		RECT	14.965 79.535 15.015 79.665 ;
		RECT	19.485 77.115 19.535 77.245 ;
		RECT	19.485 79.535 19.535 79.665 ;
		RECT	14.565 80.225 14.615 80.355 ;
		RECT	19.885 80.225 19.935 80.355 ;
		RECT	14.765 79.995 14.815 80.125 ;
		RECT	14.765 82.415 14.815 82.545 ;
		RECT	19.685 79.995 19.735 80.125 ;
		RECT	19.685 82.415 19.735 82.545 ;
		RECT	14.965 79.995 15.015 80.125 ;
		RECT	14.965 82.415 15.015 82.545 ;
		RECT	19.485 79.995 19.535 80.125 ;
		RECT	19.485 82.415 19.535 82.545 ;
		RECT	14.565 83.105 14.615 83.235 ;
		RECT	19.885 83.105 19.935 83.235 ;
		RECT	14.765 82.875 14.815 83.005 ;
		RECT	14.765 85.295 14.815 85.425 ;
		RECT	19.685 82.875 19.735 83.005 ;
		RECT	19.685 85.295 19.735 85.425 ;
		RECT	14.965 82.875 15.015 83.005 ;
		RECT	14.965 85.295 15.015 85.425 ;
		RECT	19.485 82.875 19.535 83.005 ;
		RECT	19.485 85.295 19.535 85.425 ;
		RECT	14.565 85.985 14.615 86.115 ;
		RECT	19.885 85.985 19.935 86.115 ;
		RECT	14.765 85.755 14.815 85.885 ;
		RECT	14.765 88.175 14.815 88.305 ;
		RECT	19.685 85.755 19.735 85.885 ;
		RECT	19.685 88.175 19.735 88.305 ;
		RECT	14.965 85.755 15.015 85.885 ;
		RECT	14.965 88.175 15.015 88.305 ;
		RECT	19.485 85.755 19.535 85.885 ;
		RECT	19.485 88.175 19.535 88.305 ;
		RECT	14.565 88.865 14.615 88.995 ;
		RECT	19.885 88.865 19.935 88.995 ;
		RECT	14.765 88.635 14.815 88.765 ;
		RECT	14.765 91.055 14.815 91.185 ;
		RECT	19.685 88.635 19.735 88.765 ;
		RECT	19.685 91.055 19.735 91.185 ;
		RECT	14.965 88.635 15.015 88.765 ;
		RECT	14.965 91.055 15.015 91.185 ;
		RECT	19.485 88.635 19.535 88.765 ;
		RECT	19.485 91.055 19.535 91.185 ;
		RECT	14.565 91.745 14.615 91.875 ;
		RECT	19.885 91.745 19.935 91.875 ;
		RECT	14.765 91.515 14.815 91.645 ;
		RECT	14.765 93.935 14.815 94.065 ;
		RECT	19.685 91.515 19.735 91.645 ;
		RECT	19.685 93.935 19.735 94.065 ;
		RECT	14.965 91.515 15.015 91.645 ;
		RECT	14.965 93.935 15.015 94.065 ;
		RECT	19.485 91.515 19.535 91.645 ;
		RECT	19.485 93.935 19.535 94.065 ;
		RECT	14.565 94.625 14.615 94.755 ;
		RECT	19.885 94.625 19.935 94.755 ;
		RECT	14.765 94.395 14.815 94.525 ;
		RECT	14.765 96.815 14.815 96.945 ;
		RECT	19.685 94.395 19.735 94.525 ;
		RECT	19.685 96.815 19.735 96.945 ;
		RECT	14.965 94.395 15.015 94.525 ;
		RECT	14.965 96.815 15.015 96.945 ;
		RECT	19.485 94.395 19.535 94.525 ;
		RECT	19.485 96.815 19.535 96.945 ;
		RECT	20.085 74.235 20.265 74.365 ;
		RECT	20.875 74.465 21.055 74.595 ;
		RECT	20.085 76.655 20.265 76.785 ;
		RECT	20.43 76.885 20.48 77.015 ;
		RECT	20.085 77.115 20.265 77.245 ;
		RECT	20.875 77.345 21.055 77.475 ;
		RECT	20.085 79.535 20.265 79.665 ;
		RECT	20.43 79.765 20.48 79.895 ;
		RECT	20.085 79.995 20.265 80.125 ;
		RECT	20.875 80.225 21.055 80.355 ;
		RECT	20.085 82.415 20.265 82.545 ;
		RECT	20.43 82.645 20.48 82.775 ;
		RECT	20.085 82.875 20.265 83.005 ;
		RECT	20.875 83.105 21.055 83.235 ;
		RECT	20.085 85.295 20.265 85.425 ;
		RECT	20.43 85.525 20.48 85.655 ;
		RECT	20.085 85.755 20.265 85.885 ;
		RECT	20.875 85.985 21.055 86.115 ;
		RECT	20.085 88.175 20.265 88.305 ;
		RECT	20.43 88.405 20.48 88.535 ;
		RECT	20.085 88.635 20.265 88.765 ;
		RECT	20.875 88.865 21.055 88.995 ;
		RECT	20.085 91.055 20.265 91.185 ;
		RECT	20.43 91.285 20.48 91.415 ;
		RECT	20.085 91.515 20.265 91.645 ;
		RECT	20.875 91.745 21.055 91.875 ;
		RECT	20.085 93.935 20.265 94.065 ;
		RECT	20.43 94.165 20.48 94.295 ;
		RECT	20.085 94.395 20.265 94.525 ;
		RECT	20.875 94.625 21.055 94.755 ;
		RECT	20.085 96.815 20.265 96.945 ;
		RECT	20.43 97.045 20.48 97.175 ;
		RECT	20.085 97.275 20.265 97.405 ;
		RECT	20.875 97.505 21.055 97.635 ;
		RECT	20.085 99.695 20.265 99.825 ;
		RECT	20.43 99.925 20.48 100.055 ;
		RECT	20.085 71.355 20.265 71.485 ;
		RECT	20.875 71.585 21.055 71.715 ;
		RECT	20.085 73.775 20.265 73.905 ;
		RECT	20.43 74.005 20.48 74.135 ;
		RECT	6.22 20.815 6.27 20.945 ;
		RECT	7.5 20.815 7.55 20.945 ;
		RECT	9.04 20.815 9.09 20.945 ;
		RECT	9.315 20.815 9.365 20.945 ;
		RECT	9.72 20.815 9.77 20.945 ;
		RECT	11.025 20.815 11.075 20.945 ;
		RECT	12.79 20.815 12.84 20.945 ;
		RECT	6.225 18.395 6.275 18.525 ;
		RECT	7.5 18.395 7.55 18.525 ;
		RECT	9.04 18.395 9.09 18.525 ;
		RECT	9.315 18.395 9.365 18.525 ;
		RECT	11.025 18.395 11.075 18.525 ;
		RECT	12.79 18.395 12.84 18.525 ;
		RECT	7.18 18.165 7.23 18.295 ;
		RECT	14.14 18.165 14.19 18.295 ;
		RECT	8.56 20.815 8.61 20.945 ;
		RECT	10.27 20.815 10.32 20.945 ;
		RECT	8.56 18.395 8.61 18.525 ;
		RECT	10.27 18.395 10.32 18.525 ;
		RECT	6.22 17.935 6.27 18.065 ;
		RECT	7.5 17.935 7.55 18.065 ;
		RECT	9.04 17.935 9.09 18.065 ;
		RECT	9.315 17.935 9.365 18.065 ;
		RECT	9.72 17.935 9.77 18.065 ;
		RECT	11.025 17.935 11.075 18.065 ;
		RECT	12.79 17.935 12.84 18.065 ;
		RECT	6.225 15.515 6.275 15.645 ;
		RECT	7.5 15.515 7.55 15.645 ;
		RECT	9.04 15.515 9.09 15.645 ;
		RECT	9.315 15.515 9.365 15.645 ;
		RECT	11.025 15.515 11.075 15.645 ;
		RECT	12.79 15.515 12.84 15.645 ;
		RECT	7.18 15.285 7.23 15.415 ;
		RECT	14.14 15.285 14.19 15.415 ;
		RECT	8.56 17.935 8.61 18.065 ;
		RECT	10.27 17.935 10.32 18.065 ;
		RECT	8.56 15.515 8.61 15.645 ;
		RECT	10.27 15.515 10.32 15.645 ;
		RECT	6.22 15.055 6.27 15.185 ;
		RECT	7.5 15.055 7.55 15.185 ;
		RECT	9.04 15.055 9.09 15.185 ;
		RECT	9.315 15.055 9.365 15.185 ;
		RECT	9.72 15.055 9.77 15.185 ;
		RECT	11.025 15.055 11.075 15.185 ;
		RECT	12.79 15.055 12.84 15.185 ;
		RECT	6.225 12.635 6.275 12.765 ;
		RECT	7.5 12.635 7.55 12.765 ;
		RECT	9.04 12.635 9.09 12.765 ;
		RECT	9.315 12.635 9.365 12.765 ;
		RECT	11.025 12.635 11.075 12.765 ;
		RECT	12.79 12.635 12.84 12.765 ;
		RECT	7.18 12.405 7.23 12.535 ;
		RECT	14.14 12.405 14.19 12.535 ;
		RECT	8.56 15.055 8.61 15.185 ;
		RECT	10.27 15.055 10.32 15.185 ;
		RECT	8.56 12.635 8.61 12.765 ;
		RECT	10.27 12.635 10.32 12.765 ;
		RECT	6.22 12.175 6.27 12.305 ;
		RECT	7.5 12.175 7.55 12.305 ;
		RECT	9.04 12.175 9.09 12.305 ;
		RECT	9.315 12.175 9.365 12.305 ;
		RECT	9.72 12.175 9.77 12.305 ;
		RECT	11.025 12.175 11.075 12.305 ;
		RECT	12.79 12.175 12.84 12.305 ;
		RECT	6.225 9.755 6.275 9.885 ;
		RECT	7.5 9.755 7.55 9.885 ;
		RECT	9.04 9.755 9.09 9.885 ;
		RECT	9.315 9.755 9.365 9.885 ;
		RECT	11.025 9.755 11.075 9.885 ;
		RECT	12.79 9.755 12.84 9.885 ;
		RECT	7.18 9.525 7.23 9.655 ;
		RECT	14.14 9.525 14.19 9.655 ;
		RECT	8.56 12.175 8.61 12.305 ;
		RECT	10.27 12.175 10.32 12.305 ;
		RECT	8.56 9.755 8.61 9.885 ;
		RECT	10.27 9.755 10.32 9.885 ;
		RECT	6.22 9.295 6.27 9.425 ;
		RECT	7.5 9.295 7.55 9.425 ;
		RECT	9.04 9.295 9.09 9.425 ;
		RECT	9.315 9.295 9.365 9.425 ;
		RECT	9.72 9.295 9.77 9.425 ;
		RECT	11.025 9.295 11.075 9.425 ;
		RECT	12.79 9.295 12.84 9.425 ;
		RECT	6.225 6.875 6.275 7.005 ;
		RECT	7.5 6.875 7.55 7.005 ;
		RECT	9.04 6.875 9.09 7.005 ;
		RECT	9.315 6.875 9.365 7.005 ;
		RECT	11.025 6.875 11.075 7.005 ;
		RECT	12.79 6.875 12.84 7.005 ;
		RECT	7.18 6.645 7.23 6.775 ;
		RECT	14.14 6.645 14.19 6.775 ;
		RECT	8.56 9.295 8.61 9.425 ;
		RECT	10.27 9.295 10.32 9.425 ;
		RECT	8.56 6.875 8.61 7.005 ;
		RECT	10.27 6.875 10.32 7.005 ;
		RECT	6.22 6.415 6.27 6.545 ;
		RECT	7.5 6.415 7.55 6.545 ;
		RECT	9.04 6.415 9.09 6.545 ;
		RECT	9.315 6.415 9.365 6.545 ;
		RECT	9.72 6.415 9.77 6.545 ;
		RECT	11.025 6.415 11.075 6.545 ;
		RECT	12.79 6.415 12.84 6.545 ;
		RECT	6.225 3.995 6.275 4.125 ;
		RECT	7.5 3.995 7.55 4.125 ;
		RECT	9.04 3.995 9.09 4.125 ;
		RECT	9.315 3.995 9.365 4.125 ;
		RECT	11.025 3.995 11.075 4.125 ;
		RECT	12.79 3.995 12.84 4.125 ;
		RECT	7.18 3.765 7.23 3.895 ;
		RECT	14.14 3.765 14.19 3.895 ;
		RECT	8.56 6.415 8.61 6.545 ;
		RECT	10.27 6.415 10.32 6.545 ;
		RECT	8.56 3.995 8.61 4.125 ;
		RECT	10.27 3.995 10.32 4.125 ;
		RECT	6.22 3.535 6.27 3.665 ;
		RECT	7.5 3.535 7.55 3.665 ;
		RECT	9.04 3.535 9.09 3.665 ;
		RECT	9.315 3.535 9.365 3.665 ;
		RECT	9.72 3.535 9.77 3.665 ;
		RECT	11.025 3.535 11.075 3.665 ;
		RECT	12.79 3.535 12.84 3.665 ;
		RECT	6.225 1.115 6.275 1.245 ;
		RECT	7.5 1.115 7.55 1.245 ;
		RECT	9.04 1.115 9.09 1.245 ;
		RECT	9.315 1.115 9.365 1.245 ;
		RECT	11.025 1.115 11.075 1.245 ;
		RECT	12.79 1.115 12.84 1.245 ;
		RECT	7.18 0.885 7.23 1.015 ;
		RECT	14.14 0.885 14.19 1.015 ;
		RECT	8.56 3.535 8.61 3.665 ;
		RECT	10.27 3.535 10.32 3.665 ;
		RECT	8.56 1.115 8.61 1.245 ;
		RECT	10.27 1.115 10.32 1.245 ;
		RECT	6.22 26.575 6.27 26.705 ;
		RECT	7.5 26.575 7.55 26.705 ;
		RECT	9.04 26.575 9.09 26.705 ;
		RECT	9.315 26.575 9.365 26.705 ;
		RECT	9.72 26.575 9.77 26.705 ;
		RECT	11.025 26.575 11.075 26.705 ;
		RECT	12.79 26.575 12.84 26.705 ;
		RECT	6.225 24.155 6.275 24.285 ;
		RECT	7.5 24.155 7.55 24.285 ;
		RECT	9.04 24.155 9.09 24.285 ;
		RECT	9.315 24.155 9.365 24.285 ;
		RECT	11.025 24.155 11.075 24.285 ;
		RECT	12.79 24.155 12.84 24.285 ;
		RECT	7.18 23.925 7.23 24.055 ;
		RECT	14.14 23.925 14.19 24.055 ;
		RECT	8.56 26.575 8.61 26.705 ;
		RECT	10.27 26.575 10.32 26.705 ;
		RECT	8.56 24.155 8.61 24.285 ;
		RECT	10.27 24.155 10.32 24.285 ;
		RECT	6.22 23.695 6.27 23.825 ;
		RECT	7.5 23.695 7.55 23.825 ;
		RECT	9.04 23.695 9.09 23.825 ;
		RECT	9.315 23.695 9.365 23.825 ;
		RECT	9.72 23.695 9.77 23.825 ;
		RECT	11.025 23.695 11.075 23.825 ;
		RECT	12.79 23.695 12.84 23.825 ;
		RECT	6.225 21.275 6.275 21.405 ;
		RECT	7.5 21.275 7.55 21.405 ;
		RECT	9.04 21.275 9.09 21.405 ;
		RECT	9.315 21.275 9.365 21.405 ;
		RECT	11.025 21.275 11.075 21.405 ;
		RECT	12.79 21.275 12.84 21.405 ;
		RECT	7.18 21.045 7.23 21.175 ;
		RECT	14.14 21.045 14.19 21.175 ;
		RECT	8.56 23.695 8.61 23.825 ;
		RECT	10.27 23.695 10.32 23.825 ;
		RECT	8.56 21.275 8.61 21.405 ;
		RECT	10.27 21.275 10.32 21.405 ;
		RECT	14.33 23.695 14.38 23.825 ;
		RECT	6.22 23.235 6.27 23.365 ;
		RECT	7.5 23.235 7.55 23.365 ;
		RECT	9.04 23.235 9.09 23.365 ;
		RECT	9.315 23.235 9.365 23.365 ;
		RECT	9.72 23.235 9.77 23.365 ;
		RECT	11.025 23.235 11.075 23.365 ;
		RECT	12.79 23.235 12.84 23.365 ;
		RECT	14.33 21.275 14.38 21.405 ;
		RECT	5.675 21.045 5.725 21.175 ;
		RECT	6.065 21.045 6.115 21.175 ;
		RECT	6.725 21.045 6.775 21.175 ;
		RECT	8.42 21.045 8.47 21.175 ;
		RECT	8.77 21.045 8.82 21.175 ;
		RECT	11.555 21.045 11.605 21.175 ;
		RECT	11.815 21.045 11.865 21.175 ;
		RECT	12.52 21.045 12.57 21.175 ;
		RECT	13.98 21.045 14.03 21.175 ;
		RECT	14.33 20.815 14.38 20.945 ;
		RECT	6.22 20.355 6.27 20.485 ;
		RECT	7.5 20.355 7.55 20.485 ;
		RECT	9.04 20.355 9.09 20.485 ;
		RECT	9.315 20.355 9.365 20.485 ;
		RECT	9.72 20.355 9.77 20.485 ;
		RECT	11.025 20.355 11.075 20.485 ;
		RECT	12.79 20.355 12.84 20.485 ;
		RECT	14.33 18.395 14.38 18.525 ;
		RECT	5.675 18.165 5.725 18.295 ;
		RECT	6.065 18.165 6.115 18.295 ;
		RECT	6.725 18.165 6.775 18.295 ;
		RECT	8.42 18.165 8.47 18.295 ;
		RECT	8.77 18.165 8.82 18.295 ;
		RECT	11.555 18.165 11.605 18.295 ;
		RECT	11.815 18.165 11.865 18.295 ;
		RECT	12.52 18.165 12.57 18.295 ;
		RECT	13.98 18.165 14.03 18.295 ;
		RECT	14.33 17.935 14.38 18.065 ;
		RECT	6.22 17.475 6.27 17.605 ;
		RECT	7.5 17.475 7.55 17.605 ;
		RECT	9.04 17.475 9.09 17.605 ;
		RECT	9.315 17.475 9.365 17.605 ;
		RECT	9.72 17.475 9.77 17.605 ;
		RECT	11.025 17.475 11.075 17.605 ;
		RECT	12.79 17.475 12.84 17.605 ;
		RECT	14.33 15.515 14.38 15.645 ;
		RECT	5.675 15.285 5.725 15.415 ;
		RECT	6.065 15.285 6.115 15.415 ;
		RECT	6.725 15.285 6.775 15.415 ;
		RECT	8.42 15.285 8.47 15.415 ;
		RECT	8.77 15.285 8.82 15.415 ;
		RECT	11.555 15.285 11.605 15.415 ;
		RECT	11.815 15.285 11.865 15.415 ;
		RECT	12.52 15.285 12.57 15.415 ;
		RECT	13.98 15.285 14.03 15.415 ;
		RECT	14.33 15.055 14.38 15.185 ;
		RECT	6.22 14.595 6.27 14.725 ;
		RECT	7.5 14.595 7.55 14.725 ;
		RECT	9.04 14.595 9.09 14.725 ;
		RECT	9.315 14.595 9.365 14.725 ;
		RECT	9.72 14.595 9.77 14.725 ;
		RECT	11.025 14.595 11.075 14.725 ;
		RECT	12.79 14.595 12.84 14.725 ;
		RECT	14.33 12.635 14.38 12.765 ;
		RECT	5.675 12.405 5.725 12.535 ;
		RECT	6.065 12.405 6.115 12.535 ;
		RECT	6.725 12.405 6.775 12.535 ;
		RECT	8.42 12.405 8.47 12.535 ;
		RECT	8.77 12.405 8.82 12.535 ;
		RECT	11.555 12.405 11.605 12.535 ;
		RECT	11.815 12.405 11.865 12.535 ;
		RECT	12.52 12.405 12.57 12.535 ;
		RECT	13.98 12.405 14.03 12.535 ;
		RECT	14.33 12.175 14.38 12.305 ;
		RECT	6.22 11.715 6.27 11.845 ;
		RECT	7.5 11.715 7.55 11.845 ;
		RECT	9.04 11.715 9.09 11.845 ;
		RECT	9.315 11.715 9.365 11.845 ;
		RECT	9.72 11.715 9.77 11.845 ;
		RECT	11.025 11.715 11.075 11.845 ;
		RECT	12.79 11.715 12.84 11.845 ;
		RECT	14.33 9.755 14.38 9.885 ;
		RECT	5.675 9.525 5.725 9.655 ;
		RECT	6.065 9.525 6.115 9.655 ;
		RECT	6.725 9.525 6.775 9.655 ;
		RECT	8.42 9.525 8.47 9.655 ;
		RECT	8.77 9.525 8.82 9.655 ;
		RECT	11.555 9.525 11.605 9.655 ;
		RECT	11.815 9.525 11.865 9.655 ;
		RECT	12.52 9.525 12.57 9.655 ;
		RECT	13.98 9.525 14.03 9.655 ;
		RECT	14.33 9.295 14.38 9.425 ;
		RECT	6.22 8.835 6.27 8.965 ;
		RECT	7.5 8.835 7.55 8.965 ;
		RECT	9.04 8.835 9.09 8.965 ;
		RECT	9.315 8.835 9.365 8.965 ;
		RECT	9.72 8.835 9.77 8.965 ;
		RECT	11.025 8.835 11.075 8.965 ;
		RECT	12.79 8.835 12.84 8.965 ;
		RECT	14.33 6.875 14.38 7.005 ;
		RECT	5.675 6.645 5.725 6.775 ;
		RECT	6.065 6.645 6.115 6.775 ;
		RECT	6.725 6.645 6.775 6.775 ;
		RECT	8.42 6.645 8.47 6.775 ;
		RECT	8.77 6.645 8.82 6.775 ;
		RECT	11.555 6.645 11.605 6.775 ;
		RECT	11.815 6.645 11.865 6.775 ;
		RECT	12.52 6.645 12.57 6.775 ;
		RECT	13.98 6.645 14.03 6.775 ;
		RECT	14.33 6.415 14.38 6.545 ;
		RECT	6.22 5.955 6.27 6.085 ;
		RECT	7.5 5.955 7.55 6.085 ;
		RECT	9.04 5.955 9.09 6.085 ;
		RECT	9.315 5.955 9.365 6.085 ;
		RECT	9.72 5.955 9.77 6.085 ;
		RECT	11.025 5.955 11.075 6.085 ;
		RECT	12.79 5.955 12.84 6.085 ;
		RECT	14.33 3.995 14.38 4.125 ;
		RECT	5.675 3.765 5.725 3.895 ;
		RECT	6.065 3.765 6.115 3.895 ;
		RECT	6.725 3.765 6.775 3.895 ;
		RECT	8.42 3.765 8.47 3.895 ;
		RECT	8.77 3.765 8.82 3.895 ;
		RECT	11.555 3.765 11.605 3.895 ;
		RECT	11.815 3.765 11.865 3.895 ;
		RECT	12.52 3.765 12.57 3.895 ;
		RECT	13.98 3.765 14.03 3.895 ;
		RECT	14.33 3.535 14.38 3.665 ;
		RECT	6.22 3.075 6.27 3.205 ;
		RECT	7.5 3.075 7.55 3.205 ;
		RECT	9.04 3.075 9.09 3.205 ;
		RECT	9.315 3.075 9.365 3.205 ;
		RECT	9.72 3.075 9.77 3.205 ;
		RECT	11.025 3.075 11.075 3.205 ;
		RECT	12.79 3.075 12.84 3.205 ;
		RECT	14.33 1.115 14.38 1.245 ;
		RECT	5.675 0.885 5.725 1.015 ;
		RECT	6.065 0.885 6.115 1.015 ;
		RECT	6.725 0.885 6.775 1.015 ;
		RECT	8.42 0.885 8.47 1.015 ;
		RECT	8.77 0.885 8.82 1.015 ;
		RECT	11.555 0.885 11.605 1.015 ;
		RECT	11.815 0.885 11.865 1.015 ;
		RECT	12.52 0.885 12.57 1.015 ;
		RECT	13.98 0.885 14.03 1.015 ;
		RECT	14.33 26.575 14.38 26.705 ;
		RECT	6.22 26.115 6.27 26.245 ;
		RECT	7.5 26.115 7.55 26.245 ;
		RECT	9.04 26.115 9.09 26.245 ;
		RECT	9.315 26.115 9.365 26.245 ;
		RECT	9.72 26.115 9.77 26.245 ;
		RECT	11.025 26.115 11.075 26.245 ;
		RECT	12.79 26.115 12.84 26.245 ;
		RECT	14.33 24.155 14.38 24.285 ;
		RECT	5.675 23.925 5.725 24.055 ;
		RECT	6.065 23.925 6.115 24.055 ;
		RECT	6.725 23.925 6.775 24.055 ;
		RECT	8.42 23.925 8.47 24.055 ;
		RECT	8.77 23.925 8.82 24.055 ;
		RECT	11.555 23.925 11.605 24.055 ;
		RECT	11.815 23.925 11.865 24.055 ;
		RECT	12.52 23.925 12.57 24.055 ;
		RECT	13.98 23.925 14.03 24.055 ;
		RECT	13.98 0.195 14.03 0.325 ;
		RECT	1.57 0.195 1.62 0.325 ;
		RECT	2.485 0.195 2.665 0.325 ;
		RECT	3.84 0.195 3.89 0.325 ;
		RECT	7.19 0.195 7.24 0.325 ;
		RECT	14.14 0.195 14.19 0.325 ;
		RECT	13.8 0.425 13.85 0.555 ;
		RECT	8.56 0.655 8.61 0.785 ;
		RECT	10.27 0.655 10.32 0.785 ;
		RECT	0.435 0.655 0.485 0.785 ;
		RECT	0.62 0.195 0.67 0.325 ;
		RECT	3.65 0.195 3.7 0.325 ;
		RECT	2.18 0.655 2.23 0.785 ;
		RECT	0.9 21.045 0.95 21.175 ;
		RECT	0.9 18.165 0.95 18.295 ;
		RECT	0.9 15.285 0.95 15.415 ;
		RECT	0.9 12.405 0.95 12.535 ;
		RECT	0.9 9.525 0.95 9.655 ;
		RECT	0.9 6.645 0.95 6.775 ;
		RECT	0.9 3.765 0.95 3.895 ;
		RECT	0.9 0.885 0.95 1.015 ;
		RECT	0.9 23.925 0.95 24.055 ;
		RECT	3.65 23.925 3.7 24.055 ;
		RECT	3.65 21.045 3.7 21.175 ;
		RECT	3.65 18.165 3.7 18.295 ;
		RECT	3.65 15.285 3.7 15.415 ;
		RECT	3.65 12.405 3.7 12.535 ;
		RECT	3.65 9.525 3.7 9.655 ;
		RECT	3.65 6.645 3.7 6.775 ;
		RECT	3.65 3.765 3.7 3.895 ;
		RECT	3.65 0.885 3.7 1.015 ;
		RECT	2.18 26.575 2.23 26.705 ;
		RECT	2.18 24.155 2.23 24.285 ;
		RECT	2.18 23.695 2.23 23.825 ;
		RECT	2.18 21.275 2.23 21.405 ;
		RECT	2.18 20.815 2.23 20.945 ;
		RECT	2.18 18.395 2.23 18.525 ;
		RECT	2.18 17.935 2.23 18.065 ;
		RECT	2.18 15.515 2.23 15.645 ;
		RECT	2.18 15.055 2.23 15.185 ;
		RECT	2.18 12.635 2.23 12.765 ;
		RECT	2.18 12.175 2.23 12.305 ;
		RECT	2.18 9.755 2.23 9.885 ;
		RECT	2.18 9.295 2.23 9.425 ;
		RECT	2.18 6.875 2.23 7.005 ;
		RECT	2.18 6.415 2.23 6.545 ;
		RECT	2.18 3.995 2.23 4.125 ;
		RECT	2.18 3.535 2.23 3.665 ;
		RECT	2.18 1.115 2.23 1.245 ;
		RECT	3.06 23.695 3.11 23.825 ;
		RECT	1.085 23.235 1.135 23.365 ;
		RECT	1.405 23.275 1.455 23.325 ;
		RECT	4.47 23.275 4.6 23.325 ;
		RECT	3.06 21.275 3.11 21.405 ;
		RECT	1.57 21.045 1.62 21.175 ;
		RECT	2.58 21.045 2.63 21.175 ;
		RECT	3.84 21.045 3.89 21.175 ;
		RECT	5.675 21.045 5.725 21.175 ;
		RECT	3.06 20.815 3.11 20.945 ;
		RECT	1.085 20.355 1.135 20.485 ;
		RECT	1.405 20.395 1.455 20.445 ;
		RECT	4.47 20.395 4.6 20.445 ;
		RECT	3.06 18.395 3.11 18.525 ;
		RECT	1.57 18.165 1.62 18.295 ;
		RECT	2.58 18.165 2.63 18.295 ;
		RECT	3.84 18.165 3.89 18.295 ;
		RECT	5.675 18.165 5.725 18.295 ;
		RECT	3.06 17.935 3.11 18.065 ;
		RECT	1.085 17.475 1.135 17.605 ;
		RECT	1.405 17.515 1.455 17.565 ;
		RECT	4.47 17.515 4.6 17.565 ;
		RECT	3.06 15.515 3.11 15.645 ;
		RECT	1.57 15.285 1.62 15.415 ;
		RECT	2.58 15.285 2.63 15.415 ;
		RECT	3.84 15.285 3.89 15.415 ;
		RECT	5.675 15.285 5.725 15.415 ;
		RECT	3.06 15.055 3.11 15.185 ;
		RECT	1.085 14.595 1.135 14.725 ;
		RECT	1.405 14.635 1.455 14.685 ;
		RECT	4.47 14.635 4.6 14.685 ;
		RECT	3.06 12.635 3.11 12.765 ;
		RECT	1.57 12.405 1.62 12.535 ;
		RECT	2.58 12.405 2.63 12.535 ;
		RECT	3.84 12.405 3.89 12.535 ;
		RECT	5.675 12.405 5.725 12.535 ;
		RECT	3.06 12.175 3.11 12.305 ;
		RECT	1.085 11.715 1.135 11.845 ;
		RECT	1.405 11.755 1.455 11.805 ;
		RECT	4.47 11.755 4.6 11.805 ;
		RECT	3.06 9.755 3.11 9.885 ;
		RECT	1.57 9.525 1.62 9.655 ;
		RECT	2.58 9.525 2.63 9.655 ;
		RECT	3.84 9.525 3.89 9.655 ;
		RECT	5.675 9.525 5.725 9.655 ;
		RECT	3.06 9.295 3.11 9.425 ;
		RECT	1.085 8.835 1.135 8.965 ;
		RECT	1.405 8.875 1.455 8.925 ;
		RECT	4.47 8.875 4.6 8.925 ;
		RECT	3.06 6.875 3.11 7.005 ;
		RECT	1.57 6.645 1.62 6.775 ;
		RECT	2.58 6.645 2.63 6.775 ;
		RECT	3.84 6.645 3.89 6.775 ;
		RECT	5.675 6.645 5.725 6.775 ;
		RECT	3.06 6.415 3.11 6.545 ;
		RECT	1.085 5.955 1.135 6.085 ;
		RECT	1.405 5.995 1.455 6.045 ;
		RECT	4.47 5.995 4.6 6.045 ;
		RECT	3.06 3.995 3.11 4.125 ;
		RECT	1.57 3.765 1.62 3.895 ;
		RECT	2.58 3.765 2.63 3.895 ;
		RECT	3.84 3.765 3.89 3.895 ;
		RECT	5.675 3.765 5.725 3.895 ;
		RECT	3.06 3.535 3.11 3.665 ;
		RECT	1.085 3.075 1.135 3.205 ;
		RECT	1.405 3.115 1.455 3.165 ;
		RECT	4.47 3.115 4.6 3.165 ;
		RECT	3.06 1.115 3.11 1.245 ;
		RECT	1.57 0.885 1.62 1.015 ;
		RECT	2.58 0.885 2.63 1.015 ;
		RECT	3.84 0.885 3.89 1.015 ;
		RECT	5.675 0.885 5.725 1.015 ;
		RECT	3.06 26.575 3.11 26.705 ;
		RECT	1.085 26.115 1.135 26.245 ;
		RECT	1.405 26.155 1.455 26.205 ;
		RECT	4.47 26.155 4.6 26.205 ;
		RECT	3.06 24.155 3.11 24.285 ;
		RECT	1.57 23.925 1.62 24.055 ;
		RECT	2.58 23.925 2.63 24.055 ;
		RECT	3.84 23.925 3.89 24.055 ;
		RECT	5.675 23.925 5.725 24.055 ;
		RECT	0.435 26.115 0.485 26.245 ;
		RECT	0.435 26.575 0.485 26.705 ;
		RECT	0.435 24.155 0.485 24.285 ;
		RECT	0.435 23.235 0.485 23.365 ;
		RECT	0.435 23.695 0.485 23.825 ;
		RECT	0.435 21.275 0.485 21.405 ;
		RECT	0.435 20.355 0.485 20.485 ;
		RECT	0.435 20.815 0.485 20.945 ;
		RECT	0.435 18.395 0.485 18.525 ;
		RECT	0.435 17.475 0.485 17.605 ;
		RECT	0.435 17.935 0.485 18.065 ;
		RECT	0.435 15.515 0.485 15.645 ;
		RECT	0.435 14.595 0.485 14.725 ;
		RECT	0.435 15.055 0.485 15.185 ;
		RECT	0.435 12.635 0.485 12.765 ;
		RECT	0.435 11.715 0.485 11.845 ;
		RECT	0.435 12.175 0.485 12.305 ;
		RECT	0.435 9.755 0.485 9.885 ;
		RECT	0.435 8.835 0.485 8.965 ;
		RECT	0.435 9.295 0.485 9.425 ;
		RECT	0.435 6.875 0.485 7.005 ;
		RECT	0.435 5.955 0.485 6.085 ;
		RECT	0.435 6.415 0.485 6.545 ;
		RECT	0.435 3.995 0.485 4.125 ;
		RECT	0.435 3.075 0.485 3.205 ;
		RECT	0.435 3.535 0.485 3.665 ;
		RECT	0.435 1.115 0.485 1.245 ;
		RECT	6.22 71.355 6.27 71.485 ;
		RECT	7.5 71.355 7.55 71.485 ;
		RECT	9.04 71.355 9.09 71.485 ;
		RECT	9.315 71.355 9.365 71.485 ;
		RECT	9.72 71.355 9.77 71.485 ;
		RECT	11.025 71.355 11.075 71.485 ;
		RECT	12.79 71.355 12.84 71.485 ;
		RECT	6.225 73.775 6.275 73.905 ;
		RECT	7.5 73.775 7.55 73.905 ;
		RECT	9.04 73.775 9.09 73.905 ;
		RECT	9.315 73.775 9.365 73.905 ;
		RECT	11.025 73.775 11.075 73.905 ;
		RECT	12.79 73.775 12.84 73.905 ;
		RECT	7.18 74.005 7.23 74.135 ;
		RECT	14.14 74.005 14.19 74.135 ;
		RECT	8.56 71.355 8.61 71.485 ;
		RECT	10.27 71.355 10.32 71.485 ;
		RECT	8.56 73.775 8.61 73.905 ;
		RECT	10.27 73.775 10.32 73.905 ;
		RECT	6.22 74.235 6.27 74.365 ;
		RECT	7.5 74.235 7.55 74.365 ;
		RECT	9.04 74.235 9.09 74.365 ;
		RECT	9.315 74.235 9.365 74.365 ;
		RECT	9.72 74.235 9.77 74.365 ;
		RECT	11.025 74.235 11.075 74.365 ;
		RECT	12.79 74.235 12.84 74.365 ;
		RECT	6.225 76.655 6.275 76.785 ;
		RECT	7.5 76.655 7.55 76.785 ;
		RECT	9.04 76.655 9.09 76.785 ;
		RECT	9.315 76.655 9.365 76.785 ;
		RECT	11.025 76.655 11.075 76.785 ;
		RECT	12.79 76.655 12.84 76.785 ;
		RECT	7.18 76.885 7.23 77.015 ;
		RECT	14.14 76.885 14.19 77.015 ;
		RECT	8.56 74.235 8.61 74.365 ;
		RECT	10.27 74.235 10.32 74.365 ;
		RECT	8.56 76.655 8.61 76.785 ;
		RECT	10.27 76.655 10.32 76.785 ;
		RECT	6.22 77.115 6.27 77.245 ;
		RECT	7.5 77.115 7.55 77.245 ;
		RECT	9.04 77.115 9.09 77.245 ;
		RECT	9.315 77.115 9.365 77.245 ;
		RECT	9.72 77.115 9.77 77.245 ;
		RECT	11.025 77.115 11.075 77.245 ;
		RECT	12.79 77.115 12.84 77.245 ;
		RECT	6.225 79.535 6.275 79.665 ;
		RECT	7.5 79.535 7.55 79.665 ;
		RECT	9.04 79.535 9.09 79.665 ;
		RECT	9.315 79.535 9.365 79.665 ;
		RECT	11.025 79.535 11.075 79.665 ;
		RECT	12.79 79.535 12.84 79.665 ;
		RECT	7.18 79.765 7.23 79.895 ;
		RECT	14.14 79.765 14.19 79.895 ;
		RECT	8.56 77.115 8.61 77.245 ;
		RECT	10.27 77.115 10.32 77.245 ;
		RECT	8.56 79.535 8.61 79.665 ;
		RECT	10.27 79.535 10.32 79.665 ;
		RECT	6.22 79.995 6.27 80.125 ;
		RECT	7.5 79.995 7.55 80.125 ;
		RECT	9.04 79.995 9.09 80.125 ;
		RECT	9.315 79.995 9.365 80.125 ;
		RECT	9.72 79.995 9.77 80.125 ;
		RECT	11.025 79.995 11.075 80.125 ;
		RECT	12.79 79.995 12.84 80.125 ;
		RECT	6.225 82.415 6.275 82.545 ;
		RECT	7.5 82.415 7.55 82.545 ;
		RECT	9.04 82.415 9.09 82.545 ;
		RECT	9.315 82.415 9.365 82.545 ;
		RECT	11.025 82.415 11.075 82.545 ;
		RECT	12.79 82.415 12.84 82.545 ;
		RECT	7.18 82.645 7.23 82.775 ;
		RECT	14.14 82.645 14.19 82.775 ;
		RECT	8.56 79.995 8.61 80.125 ;
		RECT	10.27 79.995 10.32 80.125 ;
		RECT	8.56 82.415 8.61 82.545 ;
		RECT	10.27 82.415 10.32 82.545 ;
		RECT	6.22 82.875 6.27 83.005 ;
		RECT	7.5 82.875 7.55 83.005 ;
		RECT	9.04 82.875 9.09 83.005 ;
		RECT	9.315 82.875 9.365 83.005 ;
		RECT	9.72 82.875 9.77 83.005 ;
		RECT	11.025 82.875 11.075 83.005 ;
		RECT	12.79 82.875 12.84 83.005 ;
		RECT	6.225 85.295 6.275 85.425 ;
		RECT	7.5 85.295 7.55 85.425 ;
		RECT	9.04 85.295 9.09 85.425 ;
		RECT	9.315 85.295 9.365 85.425 ;
		RECT	11.025 85.295 11.075 85.425 ;
		RECT	12.79 85.295 12.84 85.425 ;
		RECT	7.18 85.525 7.23 85.655 ;
		RECT	14.14 85.525 14.19 85.655 ;
		RECT	8.56 82.875 8.61 83.005 ;
		RECT	10.27 82.875 10.32 83.005 ;
		RECT	8.56 85.295 8.61 85.425 ;
		RECT	10.27 85.295 10.32 85.425 ;
		RECT	6.22 85.755 6.27 85.885 ;
		RECT	7.5 85.755 7.55 85.885 ;
		RECT	9.04 85.755 9.09 85.885 ;
		RECT	9.315 85.755 9.365 85.885 ;
		RECT	9.72 85.755 9.77 85.885 ;
		RECT	11.025 85.755 11.075 85.885 ;
		RECT	12.79 85.755 12.84 85.885 ;
		RECT	6.225 88.175 6.275 88.305 ;
		RECT	7.5 88.175 7.55 88.305 ;
		RECT	9.04 88.175 9.09 88.305 ;
		RECT	9.315 88.175 9.365 88.305 ;
		RECT	11.025 88.175 11.075 88.305 ;
		RECT	12.79 88.175 12.84 88.305 ;
		RECT	7.18 88.405 7.23 88.535 ;
		RECT	14.14 88.405 14.19 88.535 ;
		RECT	8.56 85.755 8.61 85.885 ;
		RECT	10.27 85.755 10.32 85.885 ;
		RECT	8.56 88.175 8.61 88.305 ;
		RECT	10.27 88.175 10.32 88.305 ;
		RECT	6.22 88.635 6.27 88.765 ;
		RECT	7.5 88.635 7.55 88.765 ;
		RECT	9.04 88.635 9.09 88.765 ;
		RECT	9.315 88.635 9.365 88.765 ;
		RECT	9.72 88.635 9.77 88.765 ;
		RECT	11.025 88.635 11.075 88.765 ;
		RECT	12.79 88.635 12.84 88.765 ;
		RECT	6.225 91.055 6.275 91.185 ;
		RECT	7.5 91.055 7.55 91.185 ;
		RECT	9.04 91.055 9.09 91.185 ;
		RECT	9.315 91.055 9.365 91.185 ;
		RECT	11.025 91.055 11.075 91.185 ;
		RECT	12.79 91.055 12.84 91.185 ;
		RECT	7.18 91.285 7.23 91.415 ;
		RECT	14.14 91.285 14.19 91.415 ;
		RECT	8.56 88.635 8.61 88.765 ;
		RECT	10.27 88.635 10.32 88.765 ;
		RECT	8.56 91.055 8.61 91.185 ;
		RECT	10.27 91.055 10.32 91.185 ;
		RECT	6.22 91.515 6.27 91.645 ;
		RECT	7.5 91.515 7.55 91.645 ;
		RECT	9.04 91.515 9.09 91.645 ;
		RECT	9.315 91.515 9.365 91.645 ;
		RECT	9.72 91.515 9.77 91.645 ;
		RECT	11.025 91.515 11.075 91.645 ;
		RECT	12.79 91.515 12.84 91.645 ;
		RECT	6.225 93.935 6.275 94.065 ;
		RECT	7.5 93.935 7.55 94.065 ;
		RECT	9.04 93.935 9.09 94.065 ;
		RECT	9.315 93.935 9.365 94.065 ;
		RECT	11.025 93.935 11.075 94.065 ;
		RECT	12.79 93.935 12.84 94.065 ;
		RECT	7.18 94.165 7.23 94.295 ;
		RECT	14.14 94.165 14.19 94.295 ;
		RECT	8.56 91.515 8.61 91.645 ;
		RECT	10.27 91.515 10.32 91.645 ;
		RECT	8.56 93.935 8.61 94.065 ;
		RECT	10.27 93.935 10.32 94.065 ;
		RECT	6.22 94.395 6.27 94.525 ;
		RECT	7.5 94.395 7.55 94.525 ;
		RECT	9.04 94.395 9.09 94.525 ;
		RECT	9.315 94.395 9.365 94.525 ;
		RECT	9.72 94.395 9.77 94.525 ;
		RECT	11.025 94.395 11.075 94.525 ;
		RECT	12.79 94.395 12.84 94.525 ;
		RECT	6.225 96.815 6.275 96.945 ;
		RECT	7.5 96.815 7.55 96.945 ;
		RECT	9.04 96.815 9.09 96.945 ;
		RECT	9.315 96.815 9.365 96.945 ;
		RECT	11.025 96.815 11.075 96.945 ;
		RECT	12.79 96.815 12.84 96.945 ;
		RECT	7.18 97.045 7.23 97.175 ;
		RECT	14.14 97.045 14.19 97.175 ;
		RECT	8.56 94.395 8.61 94.525 ;
		RECT	10.27 94.395 10.32 94.525 ;
		RECT	8.56 96.815 8.61 96.945 ;
		RECT	10.27 96.815 10.32 96.945 ;
		RECT	6.22 97.275 6.27 97.405 ;
		RECT	7.5 97.275 7.55 97.405 ;
		RECT	9.04 97.275 9.09 97.405 ;
		RECT	9.315 97.275 9.365 97.405 ;
		RECT	9.72 97.275 9.77 97.405 ;
		RECT	11.025 97.275 11.075 97.405 ;
		RECT	12.79 97.275 12.84 97.405 ;
		RECT	6.225 99.695 6.275 99.825 ;
		RECT	7.5 99.695 7.55 99.825 ;
		RECT	9.04 99.695 9.09 99.825 ;
		RECT	9.315 99.695 9.365 99.825 ;
		RECT	11.025 99.695 11.075 99.825 ;
		RECT	12.79 99.695 12.84 99.825 ;
		RECT	7.18 99.925 7.23 100.055 ;
		RECT	14.14 99.925 14.19 100.055 ;
		RECT	8.56 97.275 8.61 97.405 ;
		RECT	10.27 97.275 10.32 97.405 ;
		RECT	8.56 99.695 8.61 99.825 ;
		RECT	10.27 99.695 10.32 99.825 ;
		RECT	14.33 74.235 14.38 74.365 ;
		RECT	6.22 74.695 6.27 74.825 ;
		RECT	7.5 74.695 7.55 74.825 ;
		RECT	9.04 74.695 9.09 74.825 ;
		RECT	9.315 74.695 9.365 74.825 ;
		RECT	9.72 74.695 9.77 74.825 ;
		RECT	11.025 74.695 11.075 74.825 ;
		RECT	12.79 74.695 12.84 74.825 ;
		RECT	14.33 76.655 14.38 76.785 ;
		RECT	5.675 76.885 5.725 77.015 ;
		RECT	6.065 76.885 6.115 77.015 ;
		RECT	6.725 76.885 6.775 77.015 ;
		RECT	8.42 76.885 8.47 77.015 ;
		RECT	8.77 76.885 8.82 77.015 ;
		RECT	11.555 76.885 11.605 77.015 ;
		RECT	11.815 76.885 11.865 77.015 ;
		RECT	12.52 76.885 12.57 77.015 ;
		RECT	13.98 76.885 14.03 77.015 ;
		RECT	14.33 77.115 14.38 77.245 ;
		RECT	6.22 77.575 6.27 77.705 ;
		RECT	7.5 77.575 7.55 77.705 ;
		RECT	9.04 77.575 9.09 77.705 ;
		RECT	9.315 77.575 9.365 77.705 ;
		RECT	9.72 77.575 9.77 77.705 ;
		RECT	11.025 77.575 11.075 77.705 ;
		RECT	12.79 77.575 12.84 77.705 ;
		RECT	14.33 79.535 14.38 79.665 ;
		RECT	5.675 79.765 5.725 79.895 ;
		RECT	6.065 79.765 6.115 79.895 ;
		RECT	6.725 79.765 6.775 79.895 ;
		RECT	8.42 79.765 8.47 79.895 ;
		RECT	8.77 79.765 8.82 79.895 ;
		RECT	11.555 79.765 11.605 79.895 ;
		RECT	11.815 79.765 11.865 79.895 ;
		RECT	12.52 79.765 12.57 79.895 ;
		RECT	13.98 79.765 14.03 79.895 ;
		RECT	14.33 79.995 14.38 80.125 ;
		RECT	6.22 80.455 6.27 80.585 ;
		RECT	7.5 80.455 7.55 80.585 ;
		RECT	9.04 80.455 9.09 80.585 ;
		RECT	9.315 80.455 9.365 80.585 ;
		RECT	9.72 80.455 9.77 80.585 ;
		RECT	11.025 80.455 11.075 80.585 ;
		RECT	12.79 80.455 12.84 80.585 ;
		RECT	14.33 82.415 14.38 82.545 ;
		RECT	5.675 82.645 5.725 82.775 ;
		RECT	6.065 82.645 6.115 82.775 ;
		RECT	6.725 82.645 6.775 82.775 ;
		RECT	8.42 82.645 8.47 82.775 ;
		RECT	8.77 82.645 8.82 82.775 ;
		RECT	11.555 82.645 11.605 82.775 ;
		RECT	11.815 82.645 11.865 82.775 ;
		RECT	12.52 82.645 12.57 82.775 ;
		RECT	13.98 82.645 14.03 82.775 ;
		RECT	14.33 82.875 14.38 83.005 ;
		RECT	6.22 83.335 6.27 83.465 ;
		RECT	7.5 83.335 7.55 83.465 ;
		RECT	9.04 83.335 9.09 83.465 ;
		RECT	9.315 83.335 9.365 83.465 ;
		RECT	9.72 83.335 9.77 83.465 ;
		RECT	11.025 83.335 11.075 83.465 ;
		RECT	12.79 83.335 12.84 83.465 ;
		RECT	14.33 85.295 14.38 85.425 ;
		RECT	5.675 85.525 5.725 85.655 ;
		RECT	6.065 85.525 6.115 85.655 ;
		RECT	6.725 85.525 6.775 85.655 ;
		RECT	8.42 85.525 8.47 85.655 ;
		RECT	8.77 85.525 8.82 85.655 ;
		RECT	11.555 85.525 11.605 85.655 ;
		RECT	11.815 85.525 11.865 85.655 ;
		RECT	12.52 85.525 12.57 85.655 ;
		RECT	13.98 85.525 14.03 85.655 ;
		RECT	14.33 85.755 14.38 85.885 ;
		RECT	6.22 86.215 6.27 86.345 ;
		RECT	7.5 86.215 7.55 86.345 ;
		RECT	9.04 86.215 9.09 86.345 ;
		RECT	9.315 86.215 9.365 86.345 ;
		RECT	9.72 86.215 9.77 86.345 ;
		RECT	11.025 86.215 11.075 86.345 ;
		RECT	12.79 86.215 12.84 86.345 ;
		RECT	14.33 88.175 14.38 88.305 ;
		RECT	5.675 88.405 5.725 88.535 ;
		RECT	6.065 88.405 6.115 88.535 ;
		RECT	6.725 88.405 6.775 88.535 ;
		RECT	8.42 88.405 8.47 88.535 ;
		RECT	8.77 88.405 8.82 88.535 ;
		RECT	11.555 88.405 11.605 88.535 ;
		RECT	11.815 88.405 11.865 88.535 ;
		RECT	12.52 88.405 12.57 88.535 ;
		RECT	13.98 88.405 14.03 88.535 ;
		RECT	14.33 88.635 14.38 88.765 ;
		RECT	6.22 89.095 6.27 89.225 ;
		RECT	7.5 89.095 7.55 89.225 ;
		RECT	9.04 89.095 9.09 89.225 ;
		RECT	9.315 89.095 9.365 89.225 ;
		RECT	9.72 89.095 9.77 89.225 ;
		RECT	11.025 89.095 11.075 89.225 ;
		RECT	12.79 89.095 12.84 89.225 ;
		RECT	14.33 91.055 14.38 91.185 ;
		RECT	5.675 91.285 5.725 91.415 ;
		RECT	6.065 91.285 6.115 91.415 ;
		RECT	6.725 91.285 6.775 91.415 ;
		RECT	8.42 91.285 8.47 91.415 ;
		RECT	8.77 91.285 8.82 91.415 ;
		RECT	11.555 91.285 11.605 91.415 ;
		RECT	11.815 91.285 11.865 91.415 ;
		RECT	12.52 91.285 12.57 91.415 ;
		RECT	13.98 91.285 14.03 91.415 ;
		RECT	14.33 91.515 14.38 91.645 ;
		RECT	6.22 91.975 6.27 92.105 ;
		RECT	7.5 91.975 7.55 92.105 ;
		RECT	9.04 91.975 9.09 92.105 ;
		RECT	9.315 91.975 9.365 92.105 ;
		RECT	9.72 91.975 9.77 92.105 ;
		RECT	11.025 91.975 11.075 92.105 ;
		RECT	12.79 91.975 12.84 92.105 ;
		RECT	14.33 93.935 14.38 94.065 ;
		RECT	5.675 94.165 5.725 94.295 ;
		RECT	6.065 94.165 6.115 94.295 ;
		RECT	6.725 94.165 6.775 94.295 ;
		RECT	8.42 94.165 8.47 94.295 ;
		RECT	8.77 94.165 8.82 94.295 ;
		RECT	11.555 94.165 11.605 94.295 ;
		RECT	11.815 94.165 11.865 94.295 ;
		RECT	12.52 94.165 12.57 94.295 ;
		RECT	13.98 94.165 14.03 94.295 ;
		RECT	14.33 94.395 14.38 94.525 ;
		RECT	6.22 94.855 6.27 94.985 ;
		RECT	7.5 94.855 7.55 94.985 ;
		RECT	9.04 94.855 9.09 94.985 ;
		RECT	9.315 94.855 9.365 94.985 ;
		RECT	9.72 94.855 9.77 94.985 ;
		RECT	11.025 94.855 11.075 94.985 ;
		RECT	12.79 94.855 12.84 94.985 ;
		RECT	14.33 96.815 14.38 96.945 ;
		RECT	5.675 97.045 5.725 97.175 ;
		RECT	6.065 97.045 6.115 97.175 ;
		RECT	6.725 97.045 6.775 97.175 ;
		RECT	8.42 97.045 8.47 97.175 ;
		RECT	8.77 97.045 8.82 97.175 ;
		RECT	11.555 97.045 11.605 97.175 ;
		RECT	11.815 97.045 11.865 97.175 ;
		RECT	12.52 97.045 12.57 97.175 ;
		RECT	13.98 97.045 14.03 97.175 ;
		RECT	14.33 97.275 14.38 97.405 ;
		RECT	6.22 97.735 6.27 97.865 ;
		RECT	7.5 97.735 7.55 97.865 ;
		RECT	9.04 97.735 9.09 97.865 ;
		RECT	9.315 97.735 9.365 97.865 ;
		RECT	9.72 97.735 9.77 97.865 ;
		RECT	11.025 97.735 11.075 97.865 ;
		RECT	12.79 97.735 12.84 97.865 ;
		RECT	14.33 99.695 14.38 99.825 ;
		RECT	5.675 99.925 5.725 100.055 ;
		RECT	6.065 99.925 6.115 100.055 ;
		RECT	6.725 99.925 6.775 100.055 ;
		RECT	8.42 99.925 8.47 100.055 ;
		RECT	8.77 99.925 8.82 100.055 ;
		RECT	11.555 99.925 11.605 100.055 ;
		RECT	11.815 99.925 11.865 100.055 ;
		RECT	12.52 99.925 12.57 100.055 ;
		RECT	13.98 99.925 14.03 100.055 ;
		RECT	14.33 71.355 14.38 71.485 ;
		RECT	6.22 71.815 6.27 71.945 ;
		RECT	7.5 71.815 7.55 71.945 ;
		RECT	9.04 71.815 9.09 71.945 ;
		RECT	9.315 71.815 9.365 71.945 ;
		RECT	9.72 71.815 9.77 71.945 ;
		RECT	11.025 71.815 11.075 71.945 ;
		RECT	12.79 71.815 12.84 71.945 ;
		RECT	14.33 73.775 14.38 73.905 ;
		RECT	5.675 74.005 5.725 74.135 ;
		RECT	6.065 74.005 6.115 74.135 ;
		RECT	6.725 74.005 6.775 74.135 ;
		RECT	8.42 74.005 8.47 74.135 ;
		RECT	8.77 74.005 8.82 74.135 ;
		RECT	11.555 74.005 11.605 74.135 ;
		RECT	11.815 74.005 11.865 74.135 ;
		RECT	12.52 74.005 12.57 74.135 ;
		RECT	13.98 74.005 14.03 74.135 ;
		RECT	13.98 100.615 14.03 100.745 ;
		RECT	1.57 100.615 1.62 100.745 ;
		RECT	2.485 100.615 2.665 100.745 ;
		RECT	3.84 100.615 3.89 100.745 ;
		RECT	7.19 100.615 7.24 100.745 ;
		RECT	14.14 100.615 14.19 100.745 ;
		RECT	13.8 100.385 13.85 100.515 ;
		RECT	8.56 100.155 8.61 100.285 ;
		RECT	10.27 100.155 10.32 100.285 ;
		RECT	0.435 100.155 0.485 100.285 ;
		RECT	0.62 100.615 0.67 100.745 ;
		RECT	3.65 100.615 3.7 100.745 ;
		RECT	2.18 100.155 2.23 100.285 ;
		RECT	0.9 76.885 0.95 77.015 ;
		RECT	0.9 79.765 0.95 79.895 ;
		RECT	0.9 82.645 0.95 82.775 ;
		RECT	0.9 85.525 0.95 85.655 ;
		RECT	0.9 88.405 0.95 88.535 ;
		RECT	0.9 91.285 0.95 91.415 ;
		RECT	0.9 94.165 0.95 94.295 ;
		RECT	0.9 97.045 0.95 97.175 ;
		RECT	0.9 99.925 0.95 100.055 ;
		RECT	0.9 74.005 0.95 74.135 ;
		RECT	3.65 74.005 3.7 74.135 ;
		RECT	3.65 76.885 3.7 77.015 ;
		RECT	3.65 79.765 3.7 79.895 ;
		RECT	3.65 82.645 3.7 82.775 ;
		RECT	3.65 85.525 3.7 85.655 ;
		RECT	3.65 88.405 3.7 88.535 ;
		RECT	3.65 91.285 3.7 91.415 ;
		RECT	3.65 94.165 3.7 94.295 ;
		RECT	3.65 97.045 3.7 97.175 ;
		RECT	3.65 99.925 3.7 100.055 ;
		RECT	2.18 71.355 2.23 71.485 ;
		RECT	2.18 73.775 2.23 73.905 ;
		RECT	2.18 74.235 2.23 74.365 ;
		RECT	2.18 76.655 2.23 76.785 ;
		RECT	2.18 77.115 2.23 77.245 ;
		RECT	2.18 79.535 2.23 79.665 ;
		RECT	2.18 79.995 2.23 80.125 ;
		RECT	2.18 82.415 2.23 82.545 ;
		RECT	2.18 82.875 2.23 83.005 ;
		RECT	2.18 85.295 2.23 85.425 ;
		RECT	2.18 85.755 2.23 85.885 ;
		RECT	2.18 88.175 2.23 88.305 ;
		RECT	2.18 88.635 2.23 88.765 ;
		RECT	2.18 91.055 2.23 91.185 ;
		RECT	2.18 91.515 2.23 91.645 ;
		RECT	2.18 93.935 2.23 94.065 ;
		RECT	2.18 94.395 2.23 94.525 ;
		RECT	2.18 96.815 2.23 96.945 ;
		RECT	2.18 97.275 2.23 97.405 ;
		RECT	2.18 99.695 2.23 99.825 ;
		RECT	3.06 74.235 3.11 74.365 ;
		RECT	1.085 74.695 1.135 74.825 ;
		RECT	1.405 74.735 1.455 74.785 ;
		RECT	4.47 74.735 4.6 74.785 ;
		RECT	3.06 76.655 3.11 76.785 ;
		RECT	1.57 76.885 1.62 77.015 ;
		RECT	2.58 76.885 2.63 77.015 ;
		RECT	3.84 76.885 3.89 77.015 ;
		RECT	5.675 76.885 5.725 77.015 ;
		RECT	3.06 77.115 3.11 77.245 ;
		RECT	1.085 77.575 1.135 77.705 ;
		RECT	1.405 77.615 1.455 77.665 ;
		RECT	4.47 77.615 4.6 77.665 ;
		RECT	3.06 79.535 3.11 79.665 ;
		RECT	1.57 79.765 1.62 79.895 ;
		RECT	2.58 79.765 2.63 79.895 ;
		RECT	3.84 79.765 3.89 79.895 ;
		RECT	5.675 79.765 5.725 79.895 ;
		RECT	3.06 79.995 3.11 80.125 ;
		RECT	1.085 80.455 1.135 80.585 ;
		RECT	1.405 80.495 1.455 80.545 ;
		RECT	4.47 80.495 4.6 80.545 ;
		RECT	3.06 82.415 3.11 82.545 ;
		RECT	1.57 82.645 1.62 82.775 ;
		RECT	2.58 82.645 2.63 82.775 ;
		RECT	3.84 82.645 3.89 82.775 ;
		RECT	5.675 82.645 5.725 82.775 ;
		RECT	3.06 82.875 3.11 83.005 ;
		RECT	1.085 83.335 1.135 83.465 ;
		RECT	1.405 83.375 1.455 83.425 ;
		RECT	4.47 83.375 4.6 83.425 ;
		RECT	3.06 85.295 3.11 85.425 ;
		RECT	1.57 85.525 1.62 85.655 ;
		RECT	2.58 85.525 2.63 85.655 ;
		RECT	3.84 85.525 3.89 85.655 ;
		RECT	5.675 85.525 5.725 85.655 ;
		RECT	3.06 85.755 3.11 85.885 ;
		RECT	1.085 86.215 1.135 86.345 ;
		RECT	1.405 86.255 1.455 86.305 ;
		RECT	4.47 86.255 4.6 86.305 ;
		RECT	3.06 88.175 3.11 88.305 ;
		RECT	1.57 88.405 1.62 88.535 ;
		RECT	2.58 88.405 2.63 88.535 ;
		RECT	3.84 88.405 3.89 88.535 ;
		RECT	5.675 88.405 5.725 88.535 ;
		RECT	3.06 88.635 3.11 88.765 ;
		RECT	1.085 89.095 1.135 89.225 ;
		RECT	1.405 89.135 1.455 89.185 ;
		RECT	4.47 89.135 4.6 89.185 ;
		RECT	3.06 91.055 3.11 91.185 ;
		RECT	1.57 91.285 1.62 91.415 ;
		RECT	2.58 91.285 2.63 91.415 ;
		RECT	3.84 91.285 3.89 91.415 ;
		RECT	5.675 91.285 5.725 91.415 ;
		RECT	3.06 91.515 3.11 91.645 ;
		RECT	1.085 91.975 1.135 92.105 ;
		RECT	1.405 92.015 1.455 92.065 ;
		RECT	4.47 92.015 4.6 92.065 ;
		RECT	3.06 93.935 3.11 94.065 ;
		RECT	1.57 94.165 1.62 94.295 ;
		RECT	2.58 94.165 2.63 94.295 ;
		RECT	3.84 94.165 3.89 94.295 ;
		RECT	5.675 94.165 5.725 94.295 ;
		RECT	3.06 94.395 3.11 94.525 ;
		RECT	1.085 94.855 1.135 94.985 ;
		RECT	1.405 94.895 1.455 94.945 ;
		RECT	4.47 94.895 4.6 94.945 ;
		RECT	3.06 96.815 3.11 96.945 ;
		RECT	1.57 97.045 1.62 97.175 ;
		RECT	2.58 97.045 2.63 97.175 ;
		RECT	3.84 97.045 3.89 97.175 ;
		RECT	5.675 97.045 5.725 97.175 ;
		RECT	3.06 97.275 3.11 97.405 ;
		RECT	1.085 97.735 1.135 97.865 ;
		RECT	1.405 97.775 1.455 97.825 ;
		RECT	4.47 97.775 4.6 97.825 ;
		RECT	3.06 99.695 3.11 99.825 ;
		RECT	1.57 99.925 1.62 100.055 ;
		RECT	2.58 99.925 2.63 100.055 ;
		RECT	3.84 99.925 3.89 100.055 ;
		RECT	5.675 99.925 5.725 100.055 ;
		RECT	3.06 71.355 3.11 71.485 ;
		RECT	1.085 71.815 1.135 71.945 ;
		RECT	1.405 71.855 1.455 71.905 ;
		RECT	4.47 71.855 4.6 71.905 ;
		RECT	3.06 73.775 3.11 73.905 ;
		RECT	1.57 74.005 1.62 74.135 ;
		RECT	2.58 74.005 2.63 74.135 ;
		RECT	3.84 74.005 3.89 74.135 ;
		RECT	5.675 74.005 5.725 74.135 ;
		RECT	0.435 71.815 0.485 71.945 ;
		RECT	0.435 71.355 0.485 71.485 ;
		RECT	0.435 73.775 0.485 73.905 ;
		RECT	0.435 74.695 0.485 74.825 ;
		RECT	0.435 74.235 0.485 74.365 ;
		RECT	0.435 76.655 0.485 76.785 ;
		RECT	0.435 77.575 0.485 77.705 ;
		RECT	0.435 77.115 0.485 77.245 ;
		RECT	0.435 79.535 0.485 79.665 ;
		RECT	0.435 80.455 0.485 80.585 ;
		RECT	0.435 79.995 0.485 80.125 ;
		RECT	0.435 82.415 0.485 82.545 ;
		RECT	0.435 83.335 0.485 83.465 ;
		RECT	0.435 82.875 0.485 83.005 ;
		RECT	0.435 85.295 0.485 85.425 ;
		RECT	0.435 86.215 0.485 86.345 ;
		RECT	0.435 85.755 0.485 85.885 ;
		RECT	0.435 88.175 0.485 88.305 ;
		RECT	0.435 89.095 0.485 89.225 ;
		RECT	0.435 88.635 0.485 88.765 ;
		RECT	0.435 91.055 0.485 91.185 ;
		RECT	0.435 91.975 0.485 92.105 ;
		RECT	0.435 91.515 0.485 91.645 ;
		RECT	0.435 93.935 0.485 94.065 ;
		RECT	0.435 94.855 0.485 94.985 ;
		RECT	0.435 94.395 0.485 94.525 ;
		RECT	0.435 96.815 0.485 96.945 ;
		RECT	0.435 97.735 0.485 97.865 ;
		RECT	0.435 97.275 0.485 97.405 ;
		RECT	0.435 99.695 0.485 99.825 ;
		RECT	20.085 28.475 20.265 28.605 ;
		RECT	20.08 34.46 20.21 34.64 ;
		RECT	20.08 63.49 20.21 63.67 ;
		RECT	20.085 69.455 20.265 69.585 ;
		RECT	20.395 30.055 20.575 30.185 ;
		RECT	20.53 32.06 20.58 32.19 ;
		RECT	20.53 34.975 20.58 35.105 ;
		RECT	20.53 35.96 20.58 36.09 ;
		RECT	20.53 37.93 20.58 38.06 ;
		RECT	20.53 38.91 20.58 39.04 ;
		RECT	20.53 39.895 20.58 40.025 ;
		RECT	20.53 42.85 20.58 42.98 ;
		RECT	20.53 50.23 20.58 50.36 ;
		RECT	20.53 51.21 20.58 51.34 ;
		RECT	20.53 55.15 20.58 55.28 ;
		RECT	20.53 58.1 20.58 58.23 ;
		RECT	20.53 59.085 20.58 59.215 ;
		RECT	20.53 60.07 20.58 60.2 ;
		RECT	20.53 62.035 20.58 62.165 ;
		RECT	20.53 63.02 20.58 63.15 ;
		RECT	20.53 65.94 20.58 66.07 ;
		RECT	20.395 67.94 20.575 68.07 ;
		RECT	20.875 28.705 21.055 28.835 ;
		RECT	20.875 69.225 21.055 69.355 ;
		RECT	20.085 29.18 20.265 29.31 ;
		RECT	20.11 68.72 20.24 68.9 ;
		RECT	20.12 31.515 20.17 31.645 ;
		RECT	20.12 35.47 20.17 35.6 ;
		RECT	20.12 39.405 20.17 39.535 ;
		RECT	20.12 43.34 20.17 43.47 ;
		RECT	20.12 47.275 20.17 47.405 ;
		RECT	20.12 50.72 20.17 50.85 ;
		RECT	20.12 54.655 20.17 54.785 ;
		RECT	20.12 58.595 20.17 58.725 ;
		RECT	20.12 62.53 20.17 62.66 ;
		RECT	20.12 66.48 20.17 66.61 ;
		RECT	14.965 28.475 15.015 28.605 ;
		RECT	19.485 28.475 19.535 28.605 ;
		RECT	14.765 28.475 14.815 28.605 ;
		RECT	19.685 28.475 19.735 28.605 ;
		RECT	14.965 69.455 15.015 69.585 ;
		RECT	19.485 69.455 19.535 69.585 ;
		RECT	14.765 69.455 14.815 69.585 ;
		RECT	19.685 69.455 19.735 69.585 ;
		RECT	20.395 28.245 20.575 28.375 ;
		RECT	20.7 28.705 20.75 28.835 ;
		RECT	20.085 29.565 20.265 29.695 ;
		RECT	20.9 30.34 21.03 30.39 ;
		RECT	20.085 30.545 20.265 30.675 ;
		RECT	20.39 31.04 20.44 31.17 ;
		RECT	20.9 31.32 21.03 31.37 ;
		RECT	20.685 31.79 20.735 31.92 ;
		RECT	20.335 31.79 20.385 31.92 ;
		RECT	20.12 32.515 20.17 32.645 ;
		RECT	20.875 33.01 21.055 33.14 ;
		RECT	20.12 33.5 20.17 33.63 ;
		RECT	20.08 33.785 20.21 33.835 ;
		RECT	20.875 33.99 21.055 34.12 ;
		RECT	20.12 36.455 20.17 36.585 ;
		RECT	20.875 36.945 21.055 37.075 ;
		RECT	20.12 37.435 20.17 37.565 ;
		RECT	20.12 38.42 20.17 38.55 ;
		RECT	20.12 40.39 20.17 40.52 ;
		RECT	20.875 40.88 21.055 41.01 ;
		RECT	20.12 41.37 20.17 41.5 ;
		RECT	20.875 41.865 21.055 41.995 ;
		RECT	20.12 42.355 20.17 42.485 ;
		RECT	20.53 43.835 20.58 43.965 ;
		RECT	20.12 44.33 20.17 44.46 ;
		RECT	20.875 44.815 21.055 44.945 ;
		RECT	20.12 45.31 20.17 45.44 ;
		RECT	20.505 45.785 20.555 45.915 ;
		RECT	20.685 46.095 20.735 46.225 ;
		RECT	20.335 46.095 20.385 46.225 ;
		RECT	20.345 46.41 20.395 46.54 ;
		RECT	20.9 47.07 21.03 47.12 ;
		RECT	20.9 47.565 21.03 47.615 ;
		RECT	20.12 48.26 20.17 48.39 ;
		RECT	20.875 48.75 21.055 48.88 ;
		RECT	20.875 49.245 21.055 49.375 ;
		RECT	20.12 49.735 20.17 49.865 ;
		RECT	20.9 50.515 21.03 50.565 ;
		RECT	20.9 51.005 21.03 51.055 ;
		RECT	20.345 51.525 20.395 51.655 ;
		RECT	20.685 51.87 20.735 52 ;
		RECT	20.335 51.87 20.385 52 ;
		RECT	20.12 52.685 20.17 52.815 ;
		RECT	20.875 53.18 21.055 53.31 ;
		RECT	20.12 53.675 20.17 53.805 ;
		RECT	20.53 54.165 20.58 54.295 ;
		RECT	20.12 55.64 20.17 55.77 ;
		RECT	20.875 56.135 21.055 56.265 ;
		RECT	20.12 56.625 20.17 56.755 ;
		RECT	20.875 57.115 21.055 57.245 ;
		RECT	20.12 57.61 20.17 57.74 ;
		RECT	20.12 59.575 20.17 59.705 ;
		RECT	20.12 60.56 20.17 60.69 ;
		RECT	20.875 61.055 21.055 61.185 ;
		RECT	20.12 61.545 20.17 61.675 ;
		RECT	20.08 62.32 20.21 62.37 ;
		RECT	20.08 63.8 20.21 63.85 ;
		RECT	20.875 64.005 21.055 64.135 ;
		RECT	20.08 64.29 20.21 64.34 ;
		RECT	20.12 64.495 20.17 64.625 ;
		RECT	20.875 64.955 21.055 65.085 ;
		RECT	20.12 65.48 20.17 65.61 ;
		RECT	20.685 66.21 20.735 66.34 ;
		RECT	20.335 66.21 20.385 66.34 ;
		RECT	20.9 66.755 21.03 66.805 ;
		RECT	20.39 66.955 20.44 67.085 ;
		RECT	20.085 67.45 20.265 67.58 ;
		RECT	20.9 67.735 21.03 67.785 ;
		RECT	20.085 68.435 20.265 68.565 ;
		RECT	20.7 69.225 20.75 69.355 ;
		RECT	20.395 69.685 20.575 69.815 ;
		RECT	14.965 29.18 15.015 29.31 ;
		RECT	14.99 32.515 15.04 32.645 ;
		RECT	14.99 33.5 15.04 33.63 ;
		RECT	14.99 33.785 15.04 33.835 ;
		RECT	14.99 36.455 15.04 36.585 ;
		RECT	14.99 37.435 15.04 37.565 ;
		RECT	14.99 38.42 15.04 38.55 ;
		RECT	14.99 40.39 15.04 40.52 ;
		RECT	14.99 41.37 15.04 41.5 ;
		RECT	14.99 42.355 15.04 42.485 ;
		RECT	14.99 44.33 15.04 44.46 ;
		RECT	14.99 45.31 15.04 45.44 ;
		RECT	14.965 48.26 15.015 48.39 ;
		RECT	14.965 49.735 15.015 49.865 ;
		RECT	14.99 52.685 15.04 52.815 ;
		RECT	14.99 53.675 15.04 53.805 ;
		RECT	14.99 55.64 15.04 55.77 ;
		RECT	14.99 56.625 15.04 56.755 ;
		RECT	14.99 57.61 15.04 57.74 ;
		RECT	14.99 59.575 15.04 59.705 ;
		RECT	14.99 60.56 15.04 60.69 ;
		RECT	14.99 61.545 15.04 61.675 ;
		RECT	14.99 62.32 15.04 62.37 ;
		RECT	14.99 64.495 15.04 64.625 ;
		RECT	14.99 65.48 15.04 65.61 ;
		RECT	14.965 68.745 15.015 68.875 ;
		RECT	19.485 29.18 19.535 29.31 ;
		RECT	19.465 43.315 19.595 43.495 ;
		RECT	19.465 54.63 19.595 54.81 ;
		RECT	19.465 62.505 19.595 62.685 ;
		RECT	19.485 68.745 19.535 68.875 ;
		RECT	19.875 45.785 19.925 45.915 ;
		RECT	19.875 52.21 19.925 52.34 ;
		RECT	19.7 29.565 19.75 29.695 ;
		RECT	19.7 30.545 19.75 30.675 ;
		RECT	19.7 32.515 19.75 32.645 ;
		RECT	19.7 33.5 19.75 33.63 ;
		RECT	19.7 33.785 19.75 33.835 ;
		RECT	19.7 36.455 19.75 36.585 ;
		RECT	19.7 37.435 19.75 37.565 ;
		RECT	19.7 38.42 19.75 38.55 ;
		RECT	19.7 40.39 19.75 40.52 ;
		RECT	19.7 41.37 19.75 41.5 ;
		RECT	19.7 42.355 19.75 42.485 ;
		RECT	19.7 44.33 19.75 44.46 ;
		RECT	19.7 45.31 19.75 45.44 ;
		RECT	19.7 48.26 19.75 48.39 ;
		RECT	19.7 49.735 19.75 49.865 ;
		RECT	19.7 52.685 19.75 52.815 ;
		RECT	19.7 53.675 19.75 53.805 ;
		RECT	19.7 55.64 19.75 55.77 ;
		RECT	19.7 56.625 19.75 56.755 ;
		RECT	19.7 57.61 19.75 57.74 ;
		RECT	19.7 59.575 19.75 59.705 ;
		RECT	19.7 60.56 19.75 60.69 ;
		RECT	19.7 61.545 19.75 61.675 ;
		RECT	19.7 62.32 19.75 62.37 ;
		RECT	19.465 63.49 19.595 63.67 ;
		RECT	19.7 64.495 19.75 64.625 ;
		RECT	19.7 65.48 19.75 65.61 ;
		RECT	19.7 67.45 19.75 67.58 ;
		RECT	19.7 68.435 19.75 68.565 ;
		RECT	14.765 29.565 14.815 29.695 ;
		RECT	14.765 30.545 14.815 30.675 ;
		RECT	14.74 32.515 14.79 32.645 ;
		RECT	14.74 33.5 14.79 33.63 ;
		RECT	14.74 33.785 14.79 33.835 ;
		RECT	14.74 36.455 14.79 36.585 ;
		RECT	14.74 37.435 14.79 37.565 ;
		RECT	14.74 38.42 14.79 38.55 ;
		RECT	14.74 40.39 14.79 40.52 ;
		RECT	14.74 41.37 14.79 41.5 ;
		RECT	14.74 42.355 14.79 42.485 ;
		RECT	14.74 44.33 14.79 44.46 ;
		RECT	14.74 45.31 14.79 45.44 ;
		RECT	14.765 48.26 14.815 48.39 ;
		RECT	14.765 49.735 14.815 49.865 ;
		RECT	14.74 52.685 14.79 52.815 ;
		RECT	14.74 53.675 14.79 53.805 ;
		RECT	14.74 55.64 14.79 55.77 ;
		RECT	14.74 56.625 14.79 56.755 ;
		RECT	14.74 57.61 14.79 57.74 ;
		RECT	14.74 59.575 14.79 59.705 ;
		RECT	14.74 60.56 14.79 60.69 ;
		RECT	14.74 61.545 14.79 61.675 ;
		RECT	14.74 62.32 14.79 62.37 ;
		RECT	14.74 64.495 14.79 64.625 ;
		RECT	14.74 65.48 14.79 65.61 ;
		RECT	14.765 67.45 14.815 67.58 ;
		RECT	14.765 68.435 14.815 68.565 ;
		RECT	14.565 45.785 14.615 45.915 ;
		RECT	14.565 52.21 14.615 52.34 ;
		RECT	14.965 29.565 15.015 29.695 ;
		RECT	15.335 29.565 15.385 29.695 ;
		RECT	15.875 29.565 15.925 29.695 ;
		RECT	16.415 29.565 16.465 29.695 ;
		RECT	16.955 29.565 17.005 29.695 ;
		RECT	17.495 29.565 17.545 29.695 ;
		RECT	18.035 29.565 18.085 29.695 ;
		RECT	18.575 29.565 18.625 29.695 ;
		RECT	19.115 29.565 19.165 29.695 ;
		RECT	14.565 30.34 14.615 30.39 ;
		RECT	14.965 30.545 15.015 30.675 ;
		RECT	15.335 31.04 15.385 31.17 ;
		RECT	15.875 31.04 15.925 31.17 ;
		RECT	16.415 31.04 16.465 31.17 ;
		RECT	16.955 31.04 17.005 31.17 ;
		RECT	17.495 31.04 17.545 31.17 ;
		RECT	18.035 31.04 18.085 31.17 ;
		RECT	18.575 31.04 18.625 31.17 ;
		RECT	19.115 31.04 19.165 31.17 ;
		RECT	14.565 31.32 14.615 31.37 ;
		RECT	14.99 31.515 15.04 31.645 ;
		RECT	14.865 31.79 14.915 31.92 ;
		RECT	15.335 31.79 15.385 31.92 ;
		RECT	15.875 31.79 15.925 31.92 ;
		RECT	16.415 31.79 16.465 31.92 ;
		RECT	16.955 31.79 17.005 31.92 ;
		RECT	17.495 31.79 17.545 31.92 ;
		RECT	18.035 31.79 18.085 31.92 ;
		RECT	18.575 31.79 18.625 31.92 ;
		RECT	19.115 31.79 19.165 31.92 ;
		RECT	14.565 33.01 14.615 33.14 ;
		RECT	14.565 33.99 14.615 34.12 ;
		RECT	14.745 34.485 14.795 34.615 ;
		RECT	14.99 35.47 15.04 35.6 ;
		RECT	14.565 36.945 14.615 37.075 ;
		RECT	14.99 39.405 15.04 39.535 ;
		RECT	14.565 40.855 14.615 41.035 ;
		RECT	14.565 41.84 14.615 42.025 ;
		RECT	14.99 43.315 15.04 43.495 ;
		RECT	14.565 44.79 14.615 44.97 ;
		RECT	13.8 45.785 13.85 45.915 ;
		RECT	14.865 46.095 14.915 46.225 ;
		RECT	15.335 46.095 15.385 46.225 ;
		RECT	15.875 46.095 15.925 46.225 ;
		RECT	16.415 46.095 16.465 46.225 ;
		RECT	16.955 46.095 17.005 46.225 ;
		RECT	17.495 46.095 17.545 46.225 ;
		RECT	18.035 46.095 18.085 46.225 ;
		RECT	18.575 46.095 18.625 46.225 ;
		RECT	19.115 46.095 19.165 46.225 ;
		RECT	15.335 46.41 15.385 46.54 ;
		RECT	15.875 46.41 15.925 46.54 ;
		RECT	16.415 46.41 16.465 46.54 ;
		RECT	16.955 46.41 17.005 46.54 ;
		RECT	17.495 46.41 17.545 46.54 ;
		RECT	18.035 46.41 18.085 46.54 ;
		RECT	18.575 46.41 18.625 46.54 ;
		RECT	19.115 46.41 19.165 46.54 ;
		RECT	14.565 47.07 14.615 47.12 ;
		RECT	14.965 47.275 15.015 47.405 ;
		RECT	14.565 47.565 14.615 47.615 ;
		RECT	15.335 48.26 15.385 48.39 ;
		RECT	15.875 48.26 15.925 48.39 ;
		RECT	16.415 48.26 16.465 48.39 ;
		RECT	16.955 48.26 17.005 48.39 ;
		RECT	17.495 48.26 17.545 48.39 ;
		RECT	18.035 48.26 18.085 48.39 ;
		RECT	18.575 48.26 18.625 48.39 ;
		RECT	19.115 48.26 19.165 48.39 ;
		RECT	14.565 48.72 14.615 48.91 ;
		RECT	14.565 49.215 14.615 49.405 ;
		RECT	15.335 49.735 15.385 49.865 ;
		RECT	15.875 49.735 15.925 49.865 ;
		RECT	16.415 49.735 16.465 49.865 ;
		RECT	16.955 49.735 17.005 49.865 ;
		RECT	17.495 49.735 17.545 49.865 ;
		RECT	18.035 49.735 18.085 49.865 ;
		RECT	18.575 49.735 18.625 49.865 ;
		RECT	19.115 49.735 19.165 49.865 ;
		RECT	14.565 50.515 14.615 50.565 ;
		RECT	14.965 50.72 15.015 50.85 ;
		RECT	14.565 51.005 14.615 51.055 ;
		RECT	15.335 51.525 15.385 51.655 ;
		RECT	15.875 51.525 15.925 51.655 ;
		RECT	16.415 51.525 16.465 51.655 ;
		RECT	16.955 51.525 17.005 51.655 ;
		RECT	17.495 51.525 17.545 51.655 ;
		RECT	18.035 51.525 18.085 51.655 ;
		RECT	18.575 51.525 18.625 51.655 ;
		RECT	19.115 51.525 19.165 51.655 ;
		RECT	14.865 51.87 14.915 52 ;
		RECT	15.335 51.87 15.385 52 ;
		RECT	15.875 51.87 15.925 52 ;
		RECT	16.415 51.87 16.465 52 ;
		RECT	16.955 51.87 17.005 52 ;
		RECT	17.495 51.87 17.545 52 ;
		RECT	18.035 51.87 18.085 52 ;
		RECT	18.575 51.87 18.625 52 ;
		RECT	19.115 51.87 19.165 52 ;
		RECT	13.8 52.21 13.85 52.34 ;
		RECT	14.565 53.155 14.615 53.335 ;
		RECT	14.99 54.63 15.04 54.81 ;
		RECT	14.565 56.105 14.615 56.29 ;
		RECT	14.565 57.09 14.615 57.27 ;
		RECT	14.99 58.57 15.04 58.75 ;
		RECT	14.565 61.03 14.615 61.21 ;
		RECT	14.99 62.53 15.04 62.66 ;
		RECT	14.745 63.515 14.795 63.645 ;
		RECT	14.565 64.005 14.615 64.135 ;
		RECT	14.565 64.93 14.615 65.11 ;
		RECT	14.865 66.21 14.915 66.34 ;
		RECT	15.335 66.21 15.385 66.34 ;
		RECT	15.875 66.21 15.925 66.34 ;
		RECT	16.415 66.21 16.465 66.34 ;
		RECT	16.955 66.21 17.005 66.34 ;
		RECT	17.495 66.21 17.545 66.34 ;
		RECT	18.035 66.21 18.085 66.34 ;
		RECT	18.575 66.21 18.625 66.34 ;
		RECT	19.115 66.21 19.165 66.34 ;
		RECT	14.99 66.48 15.04 66.61 ;
		RECT	14.565 66.755 14.615 66.805 ;
		RECT	15.335 66.955 15.385 67.085 ;
		RECT	15.875 66.955 15.925 67.085 ;
		RECT	16.415 66.955 16.465 67.085 ;
		RECT	16.955 66.955 17.005 67.085 ;
		RECT	17.495 66.955 17.545 67.085 ;
		RECT	18.035 66.955 18.085 67.085 ;
		RECT	18.575 66.955 18.625 67.085 ;
		RECT	19.115 66.955 19.165 67.085 ;
		RECT	14.965 67.45 15.015 67.58 ;
		RECT	14.565 67.735 14.615 67.785 ;
		RECT	14.965 68.435 15.015 68.565 ;
		RECT	15.335 68.435 15.385 68.565 ;
		RECT	15.875 68.435 15.925 68.565 ;
		RECT	16.415 68.435 16.465 68.565 ;
		RECT	16.955 68.435 17.005 68.565 ;
		RECT	17.495 68.435 17.545 68.565 ;
		RECT	18.035 68.435 18.085 68.565 ;
		RECT	18.575 68.435 18.625 68.565 ;
		RECT	19.115 68.435 19.165 68.565 ;
		RECT	19.465 29.54 19.595 29.72 ;
		RECT	19.85 30.34 19.98 30.39 ;
		RECT	19.465 30.585 19.595 30.635 ;
		RECT	19.85 31.32 19.98 31.37 ;
		RECT	19.465 32.49 19.595 32.67 ;
		RECT	19.885 33.01 19.935 33.14 ;
		RECT	19.465 33.54 19.595 33.59 ;
		RECT	19.465 33.785 19.595 33.835 ;
		RECT	19.885 33.99 19.935 34.12 ;
		RECT	19.7 34.485 19.75 34.615 ;
		RECT	19.465 36.43 19.595 36.61 ;
		RECT	19.885 36.945 19.935 37.075 ;
		RECT	19.465 37.41 19.595 37.59 ;
		RECT	19.465 38.395 19.595 38.575 ;
		RECT	19.465 40.365 19.595 40.545 ;
		RECT	19.885 40.88 19.935 41.01 ;
		RECT	19.465 41.345 19.595 41.525 ;
		RECT	19.885 41.865 19.935 41.995 ;
		RECT	19.465 42.33 19.595 42.51 ;
		RECT	19.465 44.305 19.595 44.485 ;
		RECT	19.885 44.815 19.935 44.945 ;
		RECT	19.465 45.285 19.595 45.465 ;
		RECT	19.85 47.07 19.98 47.12 ;
		RECT	19.85 47.565 19.98 47.615 ;
		RECT	19.465 48.235 19.595 48.415 ;
		RECT	19.885 48.75 19.935 48.88 ;
		RECT	19.885 49.245 19.935 49.375 ;
		RECT	19.465 49.71 19.595 49.89 ;
		RECT	19.85 50.515 19.98 50.565 ;
		RECT	19.85 51.005 19.98 51.055 ;
		RECT	19.465 52.66 19.595 52.84 ;
		RECT	19.885 53.18 19.935 53.31 ;
		RECT	19.465 53.65 19.595 53.83 ;
		RECT	19.465 55.615 19.595 55.795 ;
		RECT	19.885 56.135 19.935 56.265 ;
		RECT	19.465 56.6 19.595 56.78 ;
		RECT	19.885 57.115 19.935 57.245 ;
		RECT	19.465 57.585 19.595 57.765 ;
		RECT	19.465 59.55 19.595 59.73 ;
		RECT	19.465 60.535 19.595 60.715 ;
		RECT	19.885 61.055 19.935 61.185 ;
		RECT	19.465 61.52 19.595 61.7 ;
		RECT	19.465 62.32 19.595 62.37 ;
		RECT	19.7 63.515 19.75 63.645 ;
		RECT	19.885 64.005 19.935 64.135 ;
		RECT	19.465 64.47 19.595 64.65 ;
		RECT	19.885 64.955 19.935 65.085 ;
		RECT	19.465 65.455 19.595 65.635 ;
		RECT	19.85 66.755 19.98 66.805 ;
		RECT	19.465 67.49 19.595 67.54 ;
		RECT	19.885 67.735 19.935 67.785 ;
		RECT	19.465 68.475 19.595 68.525 ;
	END

END rf2_32x19_wm0

END LIBRARY


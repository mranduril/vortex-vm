# Copyright (c) 1993 - 2019 ARM Limited. All Rights Reserved.
# Use of this Software is subject to the terms and conditions of the
# applicable license agreement with ARM Limited.

# PhyVGen V 8.3.0
# ARM Version r4p0
# Creation Date: Thu Oct 17 15:30:20 2019


# Memory Configuration:
# ~~~~~~~~~~~~~~~~~~~~~
#  -activity_factor 50 -atf off -back_biasing off -bits 128 -bmux on
# -bus_notation on -check_instname off -diodes on -drive 6 -ema on -frequency
# 1.0 -instname rf2_32x128_wm1 -left_bus_delim "[" -mux 2 -mvt BASE -name_case
# upper -pipeline off -power_gating off -power_type otc -pwr_gnd_rename
# vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -rcols 2 -redundancy off -retention on
# -right_bus_delim "]" -rrows 0 -ser none -site_def off -top_layer m5-m10
# -words 32 -wp_size 1 -write_mask on -write_thru off -corners
# ff_0p99v_0p99v_125c,ss_0p81v_0p81v_m40c,tt_0p90v_0p90v_25c
# 

VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO rf2_32x128_wm1
	FOREIGN rf2_32x128_wm1 0 0 ;
	SYMMETRY X Y ;
	SIZE 21.165 BY 414.86 ;
	CLASS BLOCK ;
	PIN AA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 191.27 0.25 191.37 ;
			LAYER	M2 ;
			RECT	0 191.27 0.25 191.37 ;
			LAYER	M3 ;
			RECT	0 191.27 0.25 191.37 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[0]

	PIN AA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 194.3 0.25 194.4 ;
			LAYER	M2 ;
			RECT	0 194.3 0.25 194.4 ;
			LAYER	M3 ;
			RECT	0 194.3 0.25 194.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[1]

	PIN AA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 197.33 0.25 197.43 ;
			LAYER	M2 ;
			RECT	0 197.33 0.25 197.43 ;
			LAYER	M3 ;
			RECT	0 197.33 0.25 197.43 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[2]

	PIN AA[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 198.875 0.25 198.975 ;
			LAYER	M2 ;
			RECT	0 198.875 0.25 198.975 ;
			LAYER	M3 ;
			RECT	0 198.875 0.25 198.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[3]

	PIN AA[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 201.905 0.25 202.005 ;
			LAYER	M2 ;
			RECT	0 201.905 0.25 202.005 ;
			LAYER	M3 ;
			RECT	0 201.905 0.25 202.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[4]

	PIN AB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 224.185 0.25 224.285 ;
			LAYER	M2 ;
			RECT	0 224.185 0.25 224.285 ;
			LAYER	M3 ;
			RECT	0 224.185 0.25 224.285 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[0]

	PIN AB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 220.96 0.25 221.06 ;
			LAYER	M2 ;
			RECT	0 220.96 0.25 221.06 ;
			LAYER	M3 ;
			RECT	0 220.96 0.25 221.06 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[1]

	PIN AB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 218.125 0.25 218.225 ;
			LAYER	M2 ;
			RECT	0 218.125 0.25 218.225 ;
			LAYER	M3 ;
			RECT	0 218.125 0.25 218.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[2]

	PIN AB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 216.58 0.25 216.68 ;
			LAYER	M2 ;
			RECT	0 216.58 0.25 216.68 ;
			LAYER	M3 ;
			RECT	0 216.58 0.25 216.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[3]

	PIN AB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 213.55 0.25 213.65 ;
			LAYER	M2 ;
			RECT	0 213.55 0.25 213.65 ;
			LAYER	M3 ;
			RECT	0 213.55 0.25 213.65 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[4]

	PIN AYA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 191.675 0.25 191.775 ;
			LAYER	M2 ;
			RECT	0 191.675 0.25 191.775 ;
			LAYER	M3 ;
			RECT	0 191.675 0.25 191.775 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[0]

	PIN AYA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 194.705 0.25 194.805 ;
			LAYER	M2 ;
			RECT	0 194.705 0.25 194.805 ;
			LAYER	M3 ;
			RECT	0 194.705 0.25 194.805 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[1]

	PIN AYA[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 197.735 0.25 197.835 ;
			LAYER	M2 ;
			RECT	0 197.735 0.25 197.835 ;
			LAYER	M3 ;
			RECT	0 197.735 0.25 197.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[2]

	PIN AYA[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 198.5 0.25 198.6 ;
			LAYER	M2 ;
			RECT	0 198.5 0.25 198.6 ;
			LAYER	M3 ;
			RECT	0 198.5 0.25 198.6 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[3]

	PIN AYA[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 201.705 0.25 201.805 ;
			LAYER	M2 ;
			RECT	0 201.705 0.25 201.805 ;
			LAYER	M3 ;
			RECT	0 201.705 0.25 201.805 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[4]

	PIN AYB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 223.78 0.25 223.88 ;
			LAYER	M2 ;
			RECT	0 223.78 0.25 223.88 ;
			LAYER	M3 ;
			RECT	0 223.78 0.25 223.88 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[0]

	PIN AYB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 220.75 0.25 220.85 ;
			LAYER	M2 ;
			RECT	0 220.75 0.25 220.85 ;
			LAYER	M3 ;
			RECT	0 220.75 0.25 220.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[1]

	PIN AYB[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 217.75 0.25 217.85 ;
			LAYER	M2 ;
			RECT	0 217.75 0.25 217.85 ;
			LAYER	M3 ;
			RECT	0 217.75 0.25 217.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[2]

	PIN AYB[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 216.985 0.25 217.085 ;
			LAYER	M2 ;
			RECT	0 216.985 0.25 217.085 ;
			LAYER	M3 ;
			RECT	0 216.985 0.25 217.085 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[3]

	PIN AYB[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 213.925 0.25 214.025 ;
			LAYER	M2 ;
			RECT	0 213.925 0.25 214.025 ;
			LAYER	M3 ;
			RECT	0 213.925 0.25 214.025 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[4]

	PIN CENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 188.51 0.25 188.61 ;
			LAYER	M2 ;
			RECT	0 188.51 0.25 188.61 ;
			LAYER	M3 ;
			RECT	0 188.51 0.25 188.61 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENA

	PIN CENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 228.705 0.25 228.805 ;
			LAYER	M2 ;
			RECT	0 228.705 0.25 228.805 ;
			LAYER	M3 ;
			RECT	0 228.705 0.25 228.805 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENB

	PIN CENYA
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 187.1 0.25 187.2 ;
			LAYER	M2 ;
			RECT	0 187.1 0.25 187.2 ;
			LAYER	M3 ;
			RECT	0 187.1 0.25 187.2 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENYA

	PIN CENYB
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 229.25 0.25 229.35 ;
			LAYER	M2 ;
			RECT	0 229.25 0.25 229.35 ;
			LAYER	M3 ;
			RECT	0 229.25 0.25 229.35 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENYB

	PIN CLKA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 198.13 0.25 198.23 ;
			LAYER	M2 ;
			RECT	0 198.13 0.25 198.23 ;
			LAYER	M3 ;
			RECT	0 198.13 0.25 198.23 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CLKA

	PIN CLKB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 218.78 0.25 218.88 ;
			LAYER	M2 ;
			RECT	0 218.78 0.25 218.88 ;
			LAYER	M3 ;
			RECT	0 218.78 0.25 218.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CLKB

	PIN COLLDISN
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 206.3 0.25 206.4 ;
			LAYER	M2 ;
			RECT	0 206.3 0.25 206.4 ;
			LAYER	M3 ;
			RECT	0 206.3 0.25 206.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END COLLDISN

	PIN DB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 2.195 0.25 2.295 ;
			LAYER	M2 ;
			RECT	0 2.195 0.25 2.295 ;
			LAYER	M3 ;
			RECT	0 2.195 0.25 2.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[0]

	PIN DB[100]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 334.805 0.25 334.905 ;
			LAYER	M2 ;
			RECT	0 334.805 0.25 334.905 ;
			LAYER	M3 ;
			RECT	0 334.805 0.25 334.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[100]

	PIN DB[101]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 337.685 0.25 337.785 ;
			LAYER	M2 ;
			RECT	0 337.685 0.25 337.785 ;
			LAYER	M3 ;
			RECT	0 337.685 0.25 337.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[101]

	PIN DB[102]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 340.565 0.25 340.665 ;
			LAYER	M2 ;
			RECT	0 340.565 0.25 340.665 ;
			LAYER	M3 ;
			RECT	0 340.565 0.25 340.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[102]

	PIN DB[103]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 343.445 0.25 343.545 ;
			LAYER	M2 ;
			RECT	0 343.445 0.25 343.545 ;
			LAYER	M3 ;
			RECT	0 343.445 0.25 343.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[103]

	PIN DB[104]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 346.325 0.25 346.425 ;
			LAYER	M2 ;
			RECT	0 346.325 0.25 346.425 ;
			LAYER	M3 ;
			RECT	0 346.325 0.25 346.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[104]

	PIN DB[105]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 349.205 0.25 349.305 ;
			LAYER	M2 ;
			RECT	0 349.205 0.25 349.305 ;
			LAYER	M3 ;
			RECT	0 349.205 0.25 349.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[105]

	PIN DB[106]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 352.085 0.25 352.185 ;
			LAYER	M2 ;
			RECT	0 352.085 0.25 352.185 ;
			LAYER	M3 ;
			RECT	0 352.085 0.25 352.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[106]

	PIN DB[107]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 354.965 0.25 355.065 ;
			LAYER	M2 ;
			RECT	0 354.965 0.25 355.065 ;
			LAYER	M3 ;
			RECT	0 354.965 0.25 355.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[107]

	PIN DB[108]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 357.845 0.25 357.945 ;
			LAYER	M2 ;
			RECT	0 357.845 0.25 357.945 ;
			LAYER	M3 ;
			RECT	0 357.845 0.25 357.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[108]

	PIN DB[109]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 360.725 0.25 360.825 ;
			LAYER	M2 ;
			RECT	0 360.725 0.25 360.825 ;
			LAYER	M3 ;
			RECT	0 360.725 0.25 360.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[109]

	PIN DB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.995 0.25 31.095 ;
			LAYER	M2 ;
			RECT	0 30.995 0.25 31.095 ;
			LAYER	M3 ;
			RECT	0 30.995 0.25 31.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[10]

	PIN DB[110]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 363.605 0.25 363.705 ;
			LAYER	M2 ;
			RECT	0 363.605 0.25 363.705 ;
			LAYER	M3 ;
			RECT	0 363.605 0.25 363.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[110]

	PIN DB[111]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 366.485 0.25 366.585 ;
			LAYER	M2 ;
			RECT	0 366.485 0.25 366.585 ;
			LAYER	M3 ;
			RECT	0 366.485 0.25 366.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[111]

	PIN DB[112]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 369.365 0.25 369.465 ;
			LAYER	M2 ;
			RECT	0 369.365 0.25 369.465 ;
			LAYER	M3 ;
			RECT	0 369.365 0.25 369.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[112]

	PIN DB[113]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 372.245 0.25 372.345 ;
			LAYER	M2 ;
			RECT	0 372.245 0.25 372.345 ;
			LAYER	M3 ;
			RECT	0 372.245 0.25 372.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[113]

	PIN DB[114]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 375.125 0.25 375.225 ;
			LAYER	M2 ;
			RECT	0 375.125 0.25 375.225 ;
			LAYER	M3 ;
			RECT	0 375.125 0.25 375.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[114]

	PIN DB[115]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 378.005 0.25 378.105 ;
			LAYER	M2 ;
			RECT	0 378.005 0.25 378.105 ;
			LAYER	M3 ;
			RECT	0 378.005 0.25 378.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[115]

	PIN DB[116]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 380.885 0.25 380.985 ;
			LAYER	M2 ;
			RECT	0 380.885 0.25 380.985 ;
			LAYER	M3 ;
			RECT	0 380.885 0.25 380.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[116]

	PIN DB[117]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 383.765 0.25 383.865 ;
			LAYER	M2 ;
			RECT	0 383.765 0.25 383.865 ;
			LAYER	M3 ;
			RECT	0 383.765 0.25 383.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[117]

	PIN DB[118]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 386.645 0.25 386.745 ;
			LAYER	M2 ;
			RECT	0 386.645 0.25 386.745 ;
			LAYER	M3 ;
			RECT	0 386.645 0.25 386.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[118]

	PIN DB[119]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 389.525 0.25 389.625 ;
			LAYER	M2 ;
			RECT	0 389.525 0.25 389.625 ;
			LAYER	M3 ;
			RECT	0 389.525 0.25 389.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[119]

	PIN DB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.875 0.25 33.975 ;
			LAYER	M2 ;
			RECT	0 33.875 0.25 33.975 ;
			LAYER	M3 ;
			RECT	0 33.875 0.25 33.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[11]

	PIN DB[120]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 392.405 0.25 392.505 ;
			LAYER	M2 ;
			RECT	0 392.405 0.25 392.505 ;
			LAYER	M3 ;
			RECT	0 392.405 0.25 392.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[120]

	PIN DB[121]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 395.285 0.25 395.385 ;
			LAYER	M2 ;
			RECT	0 395.285 0.25 395.385 ;
			LAYER	M3 ;
			RECT	0 395.285 0.25 395.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[121]

	PIN DB[122]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 398.165 0.25 398.265 ;
			LAYER	M2 ;
			RECT	0 398.165 0.25 398.265 ;
			LAYER	M3 ;
			RECT	0 398.165 0.25 398.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[122]

	PIN DB[123]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 401.045 0.25 401.145 ;
			LAYER	M2 ;
			RECT	0 401.045 0.25 401.145 ;
			LAYER	M3 ;
			RECT	0 401.045 0.25 401.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[123]

	PIN DB[124]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 403.925 0.25 404.025 ;
			LAYER	M2 ;
			RECT	0 403.925 0.25 404.025 ;
			LAYER	M3 ;
			RECT	0 403.925 0.25 404.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[124]

	PIN DB[125]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 406.805 0.25 406.905 ;
			LAYER	M2 ;
			RECT	0 406.805 0.25 406.905 ;
			LAYER	M3 ;
			RECT	0 406.805 0.25 406.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[125]

	PIN DB[126]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 409.685 0.25 409.785 ;
			LAYER	M2 ;
			RECT	0 409.685 0.25 409.785 ;
			LAYER	M3 ;
			RECT	0 409.685 0.25 409.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[126]

	PIN DB[127]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 412.565 0.25 412.665 ;
			LAYER	M2 ;
			RECT	0 412.565 0.25 412.665 ;
			LAYER	M3 ;
			RECT	0 412.565 0.25 412.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[127]

	PIN DB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.755 0.25 36.855 ;
			LAYER	M2 ;
			RECT	0 36.755 0.25 36.855 ;
			LAYER	M3 ;
			RECT	0 36.755 0.25 36.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[12]

	PIN DB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.635 0.25 39.735 ;
			LAYER	M2 ;
			RECT	0 39.635 0.25 39.735 ;
			LAYER	M3 ;
			RECT	0 39.635 0.25 39.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[13]

	PIN DB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.515 0.25 42.615 ;
			LAYER	M2 ;
			RECT	0 42.515 0.25 42.615 ;
			LAYER	M3 ;
			RECT	0 42.515 0.25 42.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[14]

	PIN DB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 45.395 0.25 45.495 ;
			LAYER	M2 ;
			RECT	0 45.395 0.25 45.495 ;
			LAYER	M3 ;
			RECT	0 45.395 0.25 45.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[15]

	PIN DB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 48.275 0.25 48.375 ;
			LAYER	M2 ;
			RECT	0 48.275 0.25 48.375 ;
			LAYER	M3 ;
			RECT	0 48.275 0.25 48.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[16]

	PIN DB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 51.155 0.25 51.255 ;
			LAYER	M2 ;
			RECT	0 51.155 0.25 51.255 ;
			LAYER	M3 ;
			RECT	0 51.155 0.25 51.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[17]

	PIN DB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.035 0.25 54.135 ;
			LAYER	M2 ;
			RECT	0 54.035 0.25 54.135 ;
			LAYER	M3 ;
			RECT	0 54.035 0.25 54.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[18]

	PIN DB[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.915 0.25 57.015 ;
			LAYER	M2 ;
			RECT	0 56.915 0.25 57.015 ;
			LAYER	M3 ;
			RECT	0 56.915 0.25 57.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[19]

	PIN DB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 5.075 0.25 5.175 ;
			LAYER	M2 ;
			RECT	0 5.075 0.25 5.175 ;
			LAYER	M3 ;
			RECT	0 5.075 0.25 5.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[1]

	PIN DB[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.795 0.25 59.895 ;
			LAYER	M2 ;
			RECT	0 59.795 0.25 59.895 ;
			LAYER	M3 ;
			RECT	0 59.795 0.25 59.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[20]

	PIN DB[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.675 0.25 62.775 ;
			LAYER	M2 ;
			RECT	0 62.675 0.25 62.775 ;
			LAYER	M3 ;
			RECT	0 62.675 0.25 62.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[21]

	PIN DB[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.555 0.25 65.655 ;
			LAYER	M2 ;
			RECT	0 65.555 0.25 65.655 ;
			LAYER	M3 ;
			RECT	0 65.555 0.25 65.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[22]

	PIN DB[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 68.435 0.25 68.535 ;
			LAYER	M2 ;
			RECT	0 68.435 0.25 68.535 ;
			LAYER	M3 ;
			RECT	0 68.435 0.25 68.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[23]

	PIN DB[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 71.315 0.25 71.415 ;
			LAYER	M2 ;
			RECT	0 71.315 0.25 71.415 ;
			LAYER	M3 ;
			RECT	0 71.315 0.25 71.415 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[24]

	PIN DB[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 74.195 0.25 74.295 ;
			LAYER	M2 ;
			RECT	0 74.195 0.25 74.295 ;
			LAYER	M3 ;
			RECT	0 74.195 0.25 74.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[25]

	PIN DB[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 77.075 0.25 77.175 ;
			LAYER	M2 ;
			RECT	0 77.075 0.25 77.175 ;
			LAYER	M3 ;
			RECT	0 77.075 0.25 77.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[26]

	PIN DB[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.955 0.25 80.055 ;
			LAYER	M2 ;
			RECT	0 79.955 0.25 80.055 ;
			LAYER	M3 ;
			RECT	0 79.955 0.25 80.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[27]

	PIN DB[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.835 0.25 82.935 ;
			LAYER	M2 ;
			RECT	0 82.835 0.25 82.935 ;
			LAYER	M3 ;
			RECT	0 82.835 0.25 82.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[28]

	PIN DB[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 85.715 0.25 85.815 ;
			LAYER	M2 ;
			RECT	0 85.715 0.25 85.815 ;
			LAYER	M3 ;
			RECT	0 85.715 0.25 85.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[29]

	PIN DB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.955 0.25 8.055 ;
			LAYER	M2 ;
			RECT	0 7.955 0.25 8.055 ;
			LAYER	M3 ;
			RECT	0 7.955 0.25 8.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[2]

	PIN DB[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 88.595 0.25 88.695 ;
			LAYER	M2 ;
			RECT	0 88.595 0.25 88.695 ;
			LAYER	M3 ;
			RECT	0 88.595 0.25 88.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[30]

	PIN DB[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 91.475 0.25 91.575 ;
			LAYER	M2 ;
			RECT	0 91.475 0.25 91.575 ;
			LAYER	M3 ;
			RECT	0 91.475 0.25 91.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[31]

	PIN DB[32]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 94.355 0.25 94.455 ;
			LAYER	M2 ;
			RECT	0 94.355 0.25 94.455 ;
			LAYER	M3 ;
			RECT	0 94.355 0.25 94.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[32]

	PIN DB[33]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 97.235 0.25 97.335 ;
			LAYER	M2 ;
			RECT	0 97.235 0.25 97.335 ;
			LAYER	M3 ;
			RECT	0 97.235 0.25 97.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[33]

	PIN DB[34]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 100.115 0.25 100.215 ;
			LAYER	M2 ;
			RECT	0 100.115 0.25 100.215 ;
			LAYER	M3 ;
			RECT	0 100.115 0.25 100.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[34]

	PIN DB[35]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 102.995 0.25 103.095 ;
			LAYER	M2 ;
			RECT	0 102.995 0.25 103.095 ;
			LAYER	M3 ;
			RECT	0 102.995 0.25 103.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[35]

	PIN DB[36]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 105.875 0.25 105.975 ;
			LAYER	M2 ;
			RECT	0 105.875 0.25 105.975 ;
			LAYER	M3 ;
			RECT	0 105.875 0.25 105.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[36]

	PIN DB[37]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 108.755 0.25 108.855 ;
			LAYER	M2 ;
			RECT	0 108.755 0.25 108.855 ;
			LAYER	M3 ;
			RECT	0 108.755 0.25 108.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[37]

	PIN DB[38]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 111.635 0.25 111.735 ;
			LAYER	M2 ;
			RECT	0 111.635 0.25 111.735 ;
			LAYER	M3 ;
			RECT	0 111.635 0.25 111.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[38]

	PIN DB[39]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 114.515 0.25 114.615 ;
			LAYER	M2 ;
			RECT	0 114.515 0.25 114.615 ;
			LAYER	M3 ;
			RECT	0 114.515 0.25 114.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[39]

	PIN DB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.835 0.25 10.935 ;
			LAYER	M2 ;
			RECT	0 10.835 0.25 10.935 ;
			LAYER	M3 ;
			RECT	0 10.835 0.25 10.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[3]

	PIN DB[40]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 117.395 0.25 117.495 ;
			LAYER	M2 ;
			RECT	0 117.395 0.25 117.495 ;
			LAYER	M3 ;
			RECT	0 117.395 0.25 117.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[40]

	PIN DB[41]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 120.275 0.25 120.375 ;
			LAYER	M2 ;
			RECT	0 120.275 0.25 120.375 ;
			LAYER	M3 ;
			RECT	0 120.275 0.25 120.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[41]

	PIN DB[42]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 123.155 0.25 123.255 ;
			LAYER	M2 ;
			RECT	0 123.155 0.25 123.255 ;
			LAYER	M3 ;
			RECT	0 123.155 0.25 123.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[42]

	PIN DB[43]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 126.035 0.25 126.135 ;
			LAYER	M2 ;
			RECT	0 126.035 0.25 126.135 ;
			LAYER	M3 ;
			RECT	0 126.035 0.25 126.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[43]

	PIN DB[44]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 128.915 0.25 129.015 ;
			LAYER	M2 ;
			RECT	0 128.915 0.25 129.015 ;
			LAYER	M3 ;
			RECT	0 128.915 0.25 129.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[44]

	PIN DB[45]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 131.795 0.25 131.895 ;
			LAYER	M2 ;
			RECT	0 131.795 0.25 131.895 ;
			LAYER	M3 ;
			RECT	0 131.795 0.25 131.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[45]

	PIN DB[46]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 134.675 0.25 134.775 ;
			LAYER	M2 ;
			RECT	0 134.675 0.25 134.775 ;
			LAYER	M3 ;
			RECT	0 134.675 0.25 134.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[46]

	PIN DB[47]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 137.555 0.25 137.655 ;
			LAYER	M2 ;
			RECT	0 137.555 0.25 137.655 ;
			LAYER	M3 ;
			RECT	0 137.555 0.25 137.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[47]

	PIN DB[48]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 140.435 0.25 140.535 ;
			LAYER	M2 ;
			RECT	0 140.435 0.25 140.535 ;
			LAYER	M3 ;
			RECT	0 140.435 0.25 140.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[48]

	PIN DB[49]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 143.315 0.25 143.415 ;
			LAYER	M2 ;
			RECT	0 143.315 0.25 143.415 ;
			LAYER	M3 ;
			RECT	0 143.315 0.25 143.415 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[49]

	PIN DB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.715 0.25 13.815 ;
			LAYER	M2 ;
			RECT	0 13.715 0.25 13.815 ;
			LAYER	M3 ;
			RECT	0 13.715 0.25 13.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[4]

	PIN DB[50]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 146.195 0.25 146.295 ;
			LAYER	M2 ;
			RECT	0 146.195 0.25 146.295 ;
			LAYER	M3 ;
			RECT	0 146.195 0.25 146.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[50]

	PIN DB[51]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 149.075 0.25 149.175 ;
			LAYER	M2 ;
			RECT	0 149.075 0.25 149.175 ;
			LAYER	M3 ;
			RECT	0 149.075 0.25 149.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[51]

	PIN DB[52]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 151.955 0.25 152.055 ;
			LAYER	M2 ;
			RECT	0 151.955 0.25 152.055 ;
			LAYER	M3 ;
			RECT	0 151.955 0.25 152.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[52]

	PIN DB[53]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 154.835 0.25 154.935 ;
			LAYER	M2 ;
			RECT	0 154.835 0.25 154.935 ;
			LAYER	M3 ;
			RECT	0 154.835 0.25 154.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[53]

	PIN DB[54]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 157.715 0.25 157.815 ;
			LAYER	M2 ;
			RECT	0 157.715 0.25 157.815 ;
			LAYER	M3 ;
			RECT	0 157.715 0.25 157.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[54]

	PIN DB[55]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 160.595 0.25 160.695 ;
			LAYER	M2 ;
			RECT	0 160.595 0.25 160.695 ;
			LAYER	M3 ;
			RECT	0 160.595 0.25 160.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[55]

	PIN DB[56]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 163.475 0.25 163.575 ;
			LAYER	M2 ;
			RECT	0 163.475 0.25 163.575 ;
			LAYER	M3 ;
			RECT	0 163.475 0.25 163.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[56]

	PIN DB[57]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 166.355 0.25 166.455 ;
			LAYER	M2 ;
			RECT	0 166.355 0.25 166.455 ;
			LAYER	M3 ;
			RECT	0 166.355 0.25 166.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[57]

	PIN DB[58]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 169.235 0.25 169.335 ;
			LAYER	M2 ;
			RECT	0 169.235 0.25 169.335 ;
			LAYER	M3 ;
			RECT	0 169.235 0.25 169.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[58]

	PIN DB[59]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 172.115 0.25 172.215 ;
			LAYER	M2 ;
			RECT	0 172.115 0.25 172.215 ;
			LAYER	M3 ;
			RECT	0 172.115 0.25 172.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[59]

	PIN DB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.595 0.25 16.695 ;
			LAYER	M2 ;
			RECT	0 16.595 0.25 16.695 ;
			LAYER	M3 ;
			RECT	0 16.595 0.25 16.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[5]

	PIN DB[60]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 174.995 0.25 175.095 ;
			LAYER	M2 ;
			RECT	0 174.995 0.25 175.095 ;
			LAYER	M3 ;
			RECT	0 174.995 0.25 175.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[60]

	PIN DB[61]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 177.875 0.25 177.975 ;
			LAYER	M2 ;
			RECT	0 177.875 0.25 177.975 ;
			LAYER	M3 ;
			RECT	0 177.875 0.25 177.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[61]

	PIN DB[62]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 180.755 0.25 180.855 ;
			LAYER	M2 ;
			RECT	0 180.755 0.25 180.855 ;
			LAYER	M3 ;
			RECT	0 180.755 0.25 180.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[62]

	PIN DB[63]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 183.635 0.25 183.735 ;
			LAYER	M2 ;
			RECT	0 183.635 0.25 183.735 ;
			LAYER	M3 ;
			RECT	0 183.635 0.25 183.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[63]

	PIN DB[64]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 231.125 0.25 231.225 ;
			LAYER	M2 ;
			RECT	0 231.125 0.25 231.225 ;
			LAYER	M3 ;
			RECT	0 231.125 0.25 231.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[64]

	PIN DB[65]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 234.005 0.25 234.105 ;
			LAYER	M2 ;
			RECT	0 234.005 0.25 234.105 ;
			LAYER	M3 ;
			RECT	0 234.005 0.25 234.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[65]

	PIN DB[66]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 236.885 0.25 236.985 ;
			LAYER	M2 ;
			RECT	0 236.885 0.25 236.985 ;
			LAYER	M3 ;
			RECT	0 236.885 0.25 236.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[66]

	PIN DB[67]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 239.765 0.25 239.865 ;
			LAYER	M2 ;
			RECT	0 239.765 0.25 239.865 ;
			LAYER	M3 ;
			RECT	0 239.765 0.25 239.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[67]

	PIN DB[68]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 242.645 0.25 242.745 ;
			LAYER	M2 ;
			RECT	0 242.645 0.25 242.745 ;
			LAYER	M3 ;
			RECT	0 242.645 0.25 242.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[68]

	PIN DB[69]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 245.525 0.25 245.625 ;
			LAYER	M2 ;
			RECT	0 245.525 0.25 245.625 ;
			LAYER	M3 ;
			RECT	0 245.525 0.25 245.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[69]

	PIN DB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.475 0.25 19.575 ;
			LAYER	M2 ;
			RECT	0 19.475 0.25 19.575 ;
			LAYER	M3 ;
			RECT	0 19.475 0.25 19.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[6]

	PIN DB[70]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 248.405 0.25 248.505 ;
			LAYER	M2 ;
			RECT	0 248.405 0.25 248.505 ;
			LAYER	M3 ;
			RECT	0 248.405 0.25 248.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[70]

	PIN DB[71]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 251.285 0.25 251.385 ;
			LAYER	M2 ;
			RECT	0 251.285 0.25 251.385 ;
			LAYER	M3 ;
			RECT	0 251.285 0.25 251.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[71]

	PIN DB[72]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 254.165 0.25 254.265 ;
			LAYER	M2 ;
			RECT	0 254.165 0.25 254.265 ;
			LAYER	M3 ;
			RECT	0 254.165 0.25 254.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[72]

	PIN DB[73]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 257.045 0.25 257.145 ;
			LAYER	M2 ;
			RECT	0 257.045 0.25 257.145 ;
			LAYER	M3 ;
			RECT	0 257.045 0.25 257.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[73]

	PIN DB[74]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 259.925 0.25 260.025 ;
			LAYER	M2 ;
			RECT	0 259.925 0.25 260.025 ;
			LAYER	M3 ;
			RECT	0 259.925 0.25 260.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[74]

	PIN DB[75]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 262.805 0.25 262.905 ;
			LAYER	M2 ;
			RECT	0 262.805 0.25 262.905 ;
			LAYER	M3 ;
			RECT	0 262.805 0.25 262.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[75]

	PIN DB[76]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 265.685 0.25 265.785 ;
			LAYER	M2 ;
			RECT	0 265.685 0.25 265.785 ;
			LAYER	M3 ;
			RECT	0 265.685 0.25 265.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[76]

	PIN DB[77]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 268.565 0.25 268.665 ;
			LAYER	M2 ;
			RECT	0 268.565 0.25 268.665 ;
			LAYER	M3 ;
			RECT	0 268.565 0.25 268.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[77]

	PIN DB[78]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 271.445 0.25 271.545 ;
			LAYER	M2 ;
			RECT	0 271.445 0.25 271.545 ;
			LAYER	M3 ;
			RECT	0 271.445 0.25 271.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[78]

	PIN DB[79]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 274.325 0.25 274.425 ;
			LAYER	M2 ;
			RECT	0 274.325 0.25 274.425 ;
			LAYER	M3 ;
			RECT	0 274.325 0.25 274.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[79]

	PIN DB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.355 0.25 22.455 ;
			LAYER	M2 ;
			RECT	0 22.355 0.25 22.455 ;
			LAYER	M3 ;
			RECT	0 22.355 0.25 22.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[7]

	PIN DB[80]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 277.205 0.25 277.305 ;
			LAYER	M2 ;
			RECT	0 277.205 0.25 277.305 ;
			LAYER	M3 ;
			RECT	0 277.205 0.25 277.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[80]

	PIN DB[81]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 280.085 0.25 280.185 ;
			LAYER	M2 ;
			RECT	0 280.085 0.25 280.185 ;
			LAYER	M3 ;
			RECT	0 280.085 0.25 280.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[81]

	PIN DB[82]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 282.965 0.25 283.065 ;
			LAYER	M2 ;
			RECT	0 282.965 0.25 283.065 ;
			LAYER	M3 ;
			RECT	0 282.965 0.25 283.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[82]

	PIN DB[83]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 285.845 0.25 285.945 ;
			LAYER	M2 ;
			RECT	0 285.845 0.25 285.945 ;
			LAYER	M3 ;
			RECT	0 285.845 0.25 285.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[83]

	PIN DB[84]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 288.725 0.25 288.825 ;
			LAYER	M2 ;
			RECT	0 288.725 0.25 288.825 ;
			LAYER	M3 ;
			RECT	0 288.725 0.25 288.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[84]

	PIN DB[85]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 291.605 0.25 291.705 ;
			LAYER	M2 ;
			RECT	0 291.605 0.25 291.705 ;
			LAYER	M3 ;
			RECT	0 291.605 0.25 291.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[85]

	PIN DB[86]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 294.485 0.25 294.585 ;
			LAYER	M2 ;
			RECT	0 294.485 0.25 294.585 ;
			LAYER	M3 ;
			RECT	0 294.485 0.25 294.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[86]

	PIN DB[87]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 297.365 0.25 297.465 ;
			LAYER	M2 ;
			RECT	0 297.365 0.25 297.465 ;
			LAYER	M3 ;
			RECT	0 297.365 0.25 297.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[87]

	PIN DB[88]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 300.245 0.25 300.345 ;
			LAYER	M2 ;
			RECT	0 300.245 0.25 300.345 ;
			LAYER	M3 ;
			RECT	0 300.245 0.25 300.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[88]

	PIN DB[89]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 303.125 0.25 303.225 ;
			LAYER	M2 ;
			RECT	0 303.125 0.25 303.225 ;
			LAYER	M3 ;
			RECT	0 303.125 0.25 303.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[89]

	PIN DB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.235 0.25 25.335 ;
			LAYER	M2 ;
			RECT	0 25.235 0.25 25.335 ;
			LAYER	M3 ;
			RECT	0 25.235 0.25 25.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[8]

	PIN DB[90]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 306.005 0.25 306.105 ;
			LAYER	M2 ;
			RECT	0 306.005 0.25 306.105 ;
			LAYER	M3 ;
			RECT	0 306.005 0.25 306.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[90]

	PIN DB[91]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 308.885 0.25 308.985 ;
			LAYER	M2 ;
			RECT	0 308.885 0.25 308.985 ;
			LAYER	M3 ;
			RECT	0 308.885 0.25 308.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[91]

	PIN DB[92]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 311.765 0.25 311.865 ;
			LAYER	M2 ;
			RECT	0 311.765 0.25 311.865 ;
			LAYER	M3 ;
			RECT	0 311.765 0.25 311.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[92]

	PIN DB[93]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 314.645 0.25 314.745 ;
			LAYER	M2 ;
			RECT	0 314.645 0.25 314.745 ;
			LAYER	M3 ;
			RECT	0 314.645 0.25 314.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[93]

	PIN DB[94]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 317.525 0.25 317.625 ;
			LAYER	M2 ;
			RECT	0 317.525 0.25 317.625 ;
			LAYER	M3 ;
			RECT	0 317.525 0.25 317.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[94]

	PIN DB[95]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 320.405 0.25 320.505 ;
			LAYER	M2 ;
			RECT	0 320.405 0.25 320.505 ;
			LAYER	M3 ;
			RECT	0 320.405 0.25 320.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[95]

	PIN DB[96]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 323.285 0.25 323.385 ;
			LAYER	M2 ;
			RECT	0 323.285 0.25 323.385 ;
			LAYER	M3 ;
			RECT	0 323.285 0.25 323.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[96]

	PIN DB[97]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 326.165 0.25 326.265 ;
			LAYER	M2 ;
			RECT	0 326.165 0.25 326.265 ;
			LAYER	M3 ;
			RECT	0 326.165 0.25 326.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[97]

	PIN DB[98]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 329.045 0.25 329.145 ;
			LAYER	M2 ;
			RECT	0 329.045 0.25 329.145 ;
			LAYER	M3 ;
			RECT	0 329.045 0.25 329.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[98]

	PIN DB[99]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 331.925 0.25 332.025 ;
			LAYER	M2 ;
			RECT	0 331.925 0.25 332.025 ;
			LAYER	M3 ;
			RECT	0 331.925 0.25 332.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[99]

	PIN DB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 28.115 0.25 28.215 ;
			LAYER	M2 ;
			RECT	0 28.115 0.25 28.215 ;
			LAYER	M3 ;
			RECT	0 28.115 0.25 28.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[9]

	PIN DFTRAMBYP
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 225.7 0.25 225.8 ;
			LAYER	M2 ;
			RECT	0 225.7 0.25 225.8 ;
			LAYER	M3 ;
			RECT	0 225.7 0.25 225.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DFTRAMBYP

	PIN EMAA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 199.77 0.25 199.87 ;
			LAYER	M2 ;
			RECT	0 199.77 0.25 199.87 ;
			LAYER	M3 ;
			RECT	0 199.77 0.25 199.87 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[0]

	PIN EMAA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 199.57 0.25 199.67 ;
			LAYER	M2 ;
			RECT	0 199.57 0.25 199.67 ;
			LAYER	M3 ;
			RECT	0 199.57 0.25 199.67 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[1]

	PIN EMAA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 201.505 0.25 201.605 ;
			LAYER	M2 ;
			RECT	0 201.505 0.25 201.605 ;
			LAYER	M3 ;
			RECT	0 201.505 0.25 201.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[2]

	PIN EMAB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 214.305 0.25 214.405 ;
			LAYER	M2 ;
			RECT	0 214.305 0.25 214.405 ;
			LAYER	M3 ;
			RECT	0 214.305 0.25 214.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[0]

	PIN EMAB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 215.305 0.25 215.405 ;
			LAYER	M2 ;
			RECT	0 215.305 0.25 215.405 ;
			LAYER	M3 ;
			RECT	0 215.305 0.25 215.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[1]

	PIN EMAB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 212.825 0.25 212.925 ;
			LAYER	M2 ;
			RECT	0 212.825 0.25 212.925 ;
			LAYER	M3 ;
			RECT	0 212.825 0.25 212.925 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[2]

	PIN EMASA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 187.45 0.25 187.55 ;
			LAYER	M2 ;
			RECT	0 187.45 0.25 187.55 ;
			LAYER	M3 ;
			RECT	0 187.45 0.25 187.55 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMASA

	PIN QA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 2.455 0.25 2.555 ;
			LAYER	M2 ;
			RECT	0 2.455 0.25 2.555 ;
			LAYER	M3 ;
			RECT	0 2.455 0.25 2.555 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[0]

	PIN QA[100]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 334.545 0.25 334.645 ;
			LAYER	M2 ;
			RECT	0 334.545 0.25 334.645 ;
			LAYER	M3 ;
			RECT	0 334.545 0.25 334.645 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[100]

	PIN QA[101]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 337.425 0.25 337.525 ;
			LAYER	M2 ;
			RECT	0 337.425 0.25 337.525 ;
			LAYER	M3 ;
			RECT	0 337.425 0.25 337.525 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[101]

	PIN QA[102]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 340.305 0.25 340.405 ;
			LAYER	M2 ;
			RECT	0 340.305 0.25 340.405 ;
			LAYER	M3 ;
			RECT	0 340.305 0.25 340.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[102]

	PIN QA[103]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 343.185 0.25 343.285 ;
			LAYER	M2 ;
			RECT	0 343.185 0.25 343.285 ;
			LAYER	M3 ;
			RECT	0 343.185 0.25 343.285 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[103]

	PIN QA[104]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 346.065 0.25 346.165 ;
			LAYER	M2 ;
			RECT	0 346.065 0.25 346.165 ;
			LAYER	M3 ;
			RECT	0 346.065 0.25 346.165 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[104]

	PIN QA[105]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 348.945 0.25 349.045 ;
			LAYER	M2 ;
			RECT	0 348.945 0.25 349.045 ;
			LAYER	M3 ;
			RECT	0 348.945 0.25 349.045 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[105]

	PIN QA[106]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 351.825 0.25 351.925 ;
			LAYER	M2 ;
			RECT	0 351.825 0.25 351.925 ;
			LAYER	M3 ;
			RECT	0 351.825 0.25 351.925 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[106]

	PIN QA[107]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 354.705 0.25 354.805 ;
			LAYER	M2 ;
			RECT	0 354.705 0.25 354.805 ;
			LAYER	M3 ;
			RECT	0 354.705 0.25 354.805 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[107]

	PIN QA[108]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 357.585 0.25 357.685 ;
			LAYER	M2 ;
			RECT	0 357.585 0.25 357.685 ;
			LAYER	M3 ;
			RECT	0 357.585 0.25 357.685 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[108]

	PIN QA[109]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 360.465 0.25 360.565 ;
			LAYER	M2 ;
			RECT	0 360.465 0.25 360.565 ;
			LAYER	M3 ;
			RECT	0 360.465 0.25 360.565 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[109]

	PIN QA[10]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 31.255 0.25 31.355 ;
			LAYER	M2 ;
			RECT	0 31.255 0.25 31.355 ;
			LAYER	M3 ;
			RECT	0 31.255 0.25 31.355 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[10]

	PIN QA[110]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 363.345 0.25 363.445 ;
			LAYER	M2 ;
			RECT	0 363.345 0.25 363.445 ;
			LAYER	M3 ;
			RECT	0 363.345 0.25 363.445 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[110]

	PIN QA[111]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 366.225 0.25 366.325 ;
			LAYER	M2 ;
			RECT	0 366.225 0.25 366.325 ;
			LAYER	M3 ;
			RECT	0 366.225 0.25 366.325 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[111]

	PIN QA[112]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 369.105 0.25 369.205 ;
			LAYER	M2 ;
			RECT	0 369.105 0.25 369.205 ;
			LAYER	M3 ;
			RECT	0 369.105 0.25 369.205 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[112]

	PIN QA[113]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 371.985 0.25 372.085 ;
			LAYER	M2 ;
			RECT	0 371.985 0.25 372.085 ;
			LAYER	M3 ;
			RECT	0 371.985 0.25 372.085 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[113]

	PIN QA[114]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 374.865 0.25 374.965 ;
			LAYER	M2 ;
			RECT	0 374.865 0.25 374.965 ;
			LAYER	M3 ;
			RECT	0 374.865 0.25 374.965 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[114]

	PIN QA[115]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 377.745 0.25 377.845 ;
			LAYER	M2 ;
			RECT	0 377.745 0.25 377.845 ;
			LAYER	M3 ;
			RECT	0 377.745 0.25 377.845 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[115]

	PIN QA[116]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 380.625 0.25 380.725 ;
			LAYER	M2 ;
			RECT	0 380.625 0.25 380.725 ;
			LAYER	M3 ;
			RECT	0 380.625 0.25 380.725 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[116]

	PIN QA[117]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 383.505 0.25 383.605 ;
			LAYER	M2 ;
			RECT	0 383.505 0.25 383.605 ;
			LAYER	M3 ;
			RECT	0 383.505 0.25 383.605 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[117]

	PIN QA[118]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 386.385 0.25 386.485 ;
			LAYER	M2 ;
			RECT	0 386.385 0.25 386.485 ;
			LAYER	M3 ;
			RECT	0 386.385 0.25 386.485 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[118]

	PIN QA[119]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 389.265 0.25 389.365 ;
			LAYER	M2 ;
			RECT	0 389.265 0.25 389.365 ;
			LAYER	M3 ;
			RECT	0 389.265 0.25 389.365 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[119]

	PIN QA[11]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 34.135 0.25 34.235 ;
			LAYER	M2 ;
			RECT	0 34.135 0.25 34.235 ;
			LAYER	M3 ;
			RECT	0 34.135 0.25 34.235 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[11]

	PIN QA[120]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 392.145 0.25 392.245 ;
			LAYER	M2 ;
			RECT	0 392.145 0.25 392.245 ;
			LAYER	M3 ;
			RECT	0 392.145 0.25 392.245 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[120]

	PIN QA[121]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 395.025 0.25 395.125 ;
			LAYER	M2 ;
			RECT	0 395.025 0.25 395.125 ;
			LAYER	M3 ;
			RECT	0 395.025 0.25 395.125 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[121]

	PIN QA[122]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 397.905 0.25 398.005 ;
			LAYER	M2 ;
			RECT	0 397.905 0.25 398.005 ;
			LAYER	M3 ;
			RECT	0 397.905 0.25 398.005 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[122]

	PIN QA[123]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 400.785 0.25 400.885 ;
			LAYER	M2 ;
			RECT	0 400.785 0.25 400.885 ;
			LAYER	M3 ;
			RECT	0 400.785 0.25 400.885 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[123]

	PIN QA[124]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 403.665 0.25 403.765 ;
			LAYER	M2 ;
			RECT	0 403.665 0.25 403.765 ;
			LAYER	M3 ;
			RECT	0 403.665 0.25 403.765 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[124]

	PIN QA[125]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 406.545 0.25 406.645 ;
			LAYER	M2 ;
			RECT	0 406.545 0.25 406.645 ;
			LAYER	M3 ;
			RECT	0 406.545 0.25 406.645 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[125]

	PIN QA[126]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 409.425 0.25 409.525 ;
			LAYER	M2 ;
			RECT	0 409.425 0.25 409.525 ;
			LAYER	M3 ;
			RECT	0 409.425 0.25 409.525 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[126]

	PIN QA[127]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 412.305 0.25 412.405 ;
			LAYER	M2 ;
			RECT	0 412.305 0.25 412.405 ;
			LAYER	M3 ;
			RECT	0 412.305 0.25 412.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[127]

	PIN QA[12]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 37.015 0.25 37.115 ;
			LAYER	M2 ;
			RECT	0 37.015 0.25 37.115 ;
			LAYER	M3 ;
			RECT	0 37.015 0.25 37.115 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[12]

	PIN QA[13]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.895 0.25 39.995 ;
			LAYER	M2 ;
			RECT	0 39.895 0.25 39.995 ;
			LAYER	M3 ;
			RECT	0 39.895 0.25 39.995 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[13]

	PIN QA[14]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.775 0.25 42.875 ;
			LAYER	M2 ;
			RECT	0 42.775 0.25 42.875 ;
			LAYER	M3 ;
			RECT	0 42.775 0.25 42.875 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[14]

	PIN QA[15]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 45.655 0.25 45.755 ;
			LAYER	M2 ;
			RECT	0 45.655 0.25 45.755 ;
			LAYER	M3 ;
			RECT	0 45.655 0.25 45.755 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[15]

	PIN QA[16]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 48.535 0.25 48.635 ;
			LAYER	M2 ;
			RECT	0 48.535 0.25 48.635 ;
			LAYER	M3 ;
			RECT	0 48.535 0.25 48.635 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[16]

	PIN QA[17]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 51.415 0.25 51.515 ;
			LAYER	M2 ;
			RECT	0 51.415 0.25 51.515 ;
			LAYER	M3 ;
			RECT	0 51.415 0.25 51.515 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[17]

	PIN QA[18]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.295 0.25 54.395 ;
			LAYER	M2 ;
			RECT	0 54.295 0.25 54.395 ;
			LAYER	M3 ;
			RECT	0 54.295 0.25 54.395 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[18]

	PIN QA[19]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 57.175 0.25 57.275 ;
			LAYER	M2 ;
			RECT	0 57.175 0.25 57.275 ;
			LAYER	M3 ;
			RECT	0 57.175 0.25 57.275 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[19]

	PIN QA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 5.335 0.25 5.435 ;
			LAYER	M2 ;
			RECT	0 5.335 0.25 5.435 ;
			LAYER	M3 ;
			RECT	0 5.335 0.25 5.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[1]

	PIN QA[20]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.055 0.25 60.155 ;
			LAYER	M2 ;
			RECT	0 60.055 0.25 60.155 ;
			LAYER	M3 ;
			RECT	0 60.055 0.25 60.155 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[20]

	PIN QA[21]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.935 0.25 63.035 ;
			LAYER	M2 ;
			RECT	0 62.935 0.25 63.035 ;
			LAYER	M3 ;
			RECT	0 62.935 0.25 63.035 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[21]

	PIN QA[22]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.815 0.25 65.915 ;
			LAYER	M2 ;
			RECT	0 65.815 0.25 65.915 ;
			LAYER	M3 ;
			RECT	0 65.815 0.25 65.915 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[22]

	PIN QA[23]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 68.695 0.25 68.795 ;
			LAYER	M2 ;
			RECT	0 68.695 0.25 68.795 ;
			LAYER	M3 ;
			RECT	0 68.695 0.25 68.795 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[23]

	PIN QA[24]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 71.575 0.25 71.675 ;
			LAYER	M2 ;
			RECT	0 71.575 0.25 71.675 ;
			LAYER	M3 ;
			RECT	0 71.575 0.25 71.675 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[24]

	PIN QA[25]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 74.455 0.25 74.555 ;
			LAYER	M2 ;
			RECT	0 74.455 0.25 74.555 ;
			LAYER	M3 ;
			RECT	0 74.455 0.25 74.555 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[25]

	PIN QA[26]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 77.335 0.25 77.435 ;
			LAYER	M2 ;
			RECT	0 77.335 0.25 77.435 ;
			LAYER	M3 ;
			RECT	0 77.335 0.25 77.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[26]

	PIN QA[27]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 80.215 0.25 80.315 ;
			LAYER	M2 ;
			RECT	0 80.215 0.25 80.315 ;
			LAYER	M3 ;
			RECT	0 80.215 0.25 80.315 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[27]

	PIN QA[28]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 83.095 0.25 83.195 ;
			LAYER	M2 ;
			RECT	0 83.095 0.25 83.195 ;
			LAYER	M3 ;
			RECT	0 83.095 0.25 83.195 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[28]

	PIN QA[29]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 85.975 0.25 86.075 ;
			LAYER	M2 ;
			RECT	0 85.975 0.25 86.075 ;
			LAYER	M3 ;
			RECT	0 85.975 0.25 86.075 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[29]

	PIN QA[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 8.215 0.25 8.315 ;
			LAYER	M2 ;
			RECT	0 8.215 0.25 8.315 ;
			LAYER	M3 ;
			RECT	0 8.215 0.25 8.315 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[2]

	PIN QA[30]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 88.855 0.25 88.955 ;
			LAYER	M2 ;
			RECT	0 88.855 0.25 88.955 ;
			LAYER	M3 ;
			RECT	0 88.855 0.25 88.955 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[30]

	PIN QA[31]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 91.735 0.25 91.835 ;
			LAYER	M2 ;
			RECT	0 91.735 0.25 91.835 ;
			LAYER	M3 ;
			RECT	0 91.735 0.25 91.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[31]

	PIN QA[32]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 94.615 0.25 94.715 ;
			LAYER	M2 ;
			RECT	0 94.615 0.25 94.715 ;
			LAYER	M3 ;
			RECT	0 94.615 0.25 94.715 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[32]

	PIN QA[33]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 97.495 0.25 97.595 ;
			LAYER	M2 ;
			RECT	0 97.495 0.25 97.595 ;
			LAYER	M3 ;
			RECT	0 97.495 0.25 97.595 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[33]

	PIN QA[34]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 100.375 0.25 100.475 ;
			LAYER	M2 ;
			RECT	0 100.375 0.25 100.475 ;
			LAYER	M3 ;
			RECT	0 100.375 0.25 100.475 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[34]

	PIN QA[35]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 103.255 0.25 103.355 ;
			LAYER	M2 ;
			RECT	0 103.255 0.25 103.355 ;
			LAYER	M3 ;
			RECT	0 103.255 0.25 103.355 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[35]

	PIN QA[36]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 106.135 0.25 106.235 ;
			LAYER	M2 ;
			RECT	0 106.135 0.25 106.235 ;
			LAYER	M3 ;
			RECT	0 106.135 0.25 106.235 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[36]

	PIN QA[37]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 109.015 0.25 109.115 ;
			LAYER	M2 ;
			RECT	0 109.015 0.25 109.115 ;
			LAYER	M3 ;
			RECT	0 109.015 0.25 109.115 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[37]

	PIN QA[38]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 111.895 0.25 111.995 ;
			LAYER	M2 ;
			RECT	0 111.895 0.25 111.995 ;
			LAYER	M3 ;
			RECT	0 111.895 0.25 111.995 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[38]

	PIN QA[39]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 114.775 0.25 114.875 ;
			LAYER	M2 ;
			RECT	0 114.775 0.25 114.875 ;
			LAYER	M3 ;
			RECT	0 114.775 0.25 114.875 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[39]

	PIN QA[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 11.095 0.25 11.195 ;
			LAYER	M2 ;
			RECT	0 11.095 0.25 11.195 ;
			LAYER	M3 ;
			RECT	0 11.095 0.25 11.195 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[3]

	PIN QA[40]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 117.655 0.25 117.755 ;
			LAYER	M2 ;
			RECT	0 117.655 0.25 117.755 ;
			LAYER	M3 ;
			RECT	0 117.655 0.25 117.755 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[40]

	PIN QA[41]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 120.535 0.25 120.635 ;
			LAYER	M2 ;
			RECT	0 120.535 0.25 120.635 ;
			LAYER	M3 ;
			RECT	0 120.535 0.25 120.635 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[41]

	PIN QA[42]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 123.415 0.25 123.515 ;
			LAYER	M2 ;
			RECT	0 123.415 0.25 123.515 ;
			LAYER	M3 ;
			RECT	0 123.415 0.25 123.515 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[42]

	PIN QA[43]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 126.295 0.25 126.395 ;
			LAYER	M2 ;
			RECT	0 126.295 0.25 126.395 ;
			LAYER	M3 ;
			RECT	0 126.295 0.25 126.395 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[43]

	PIN QA[44]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 129.175 0.25 129.275 ;
			LAYER	M2 ;
			RECT	0 129.175 0.25 129.275 ;
			LAYER	M3 ;
			RECT	0 129.175 0.25 129.275 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[44]

	PIN QA[45]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 132.055 0.25 132.155 ;
			LAYER	M2 ;
			RECT	0 132.055 0.25 132.155 ;
			LAYER	M3 ;
			RECT	0 132.055 0.25 132.155 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[45]

	PIN QA[46]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 134.935 0.25 135.035 ;
			LAYER	M2 ;
			RECT	0 134.935 0.25 135.035 ;
			LAYER	M3 ;
			RECT	0 134.935 0.25 135.035 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[46]

	PIN QA[47]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 137.815 0.25 137.915 ;
			LAYER	M2 ;
			RECT	0 137.815 0.25 137.915 ;
			LAYER	M3 ;
			RECT	0 137.815 0.25 137.915 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[47]

	PIN QA[48]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 140.695 0.25 140.795 ;
			LAYER	M2 ;
			RECT	0 140.695 0.25 140.795 ;
			LAYER	M3 ;
			RECT	0 140.695 0.25 140.795 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[48]

	PIN QA[49]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 143.575 0.25 143.675 ;
			LAYER	M2 ;
			RECT	0 143.575 0.25 143.675 ;
			LAYER	M3 ;
			RECT	0 143.575 0.25 143.675 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[49]

	PIN QA[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.975 0.25 14.075 ;
			LAYER	M2 ;
			RECT	0 13.975 0.25 14.075 ;
			LAYER	M3 ;
			RECT	0 13.975 0.25 14.075 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[4]

	PIN QA[50]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 146.455 0.25 146.555 ;
			LAYER	M2 ;
			RECT	0 146.455 0.25 146.555 ;
			LAYER	M3 ;
			RECT	0 146.455 0.25 146.555 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[50]

	PIN QA[51]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 149.335 0.25 149.435 ;
			LAYER	M2 ;
			RECT	0 149.335 0.25 149.435 ;
			LAYER	M3 ;
			RECT	0 149.335 0.25 149.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[51]

	PIN QA[52]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 152.215 0.25 152.315 ;
			LAYER	M2 ;
			RECT	0 152.215 0.25 152.315 ;
			LAYER	M3 ;
			RECT	0 152.215 0.25 152.315 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[52]

	PIN QA[53]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 155.095 0.25 155.195 ;
			LAYER	M2 ;
			RECT	0 155.095 0.25 155.195 ;
			LAYER	M3 ;
			RECT	0 155.095 0.25 155.195 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[53]

	PIN QA[54]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 157.975 0.25 158.075 ;
			LAYER	M2 ;
			RECT	0 157.975 0.25 158.075 ;
			LAYER	M3 ;
			RECT	0 157.975 0.25 158.075 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[54]

	PIN QA[55]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 160.855 0.25 160.955 ;
			LAYER	M2 ;
			RECT	0 160.855 0.25 160.955 ;
			LAYER	M3 ;
			RECT	0 160.855 0.25 160.955 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[55]

	PIN QA[56]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 163.735 0.25 163.835 ;
			LAYER	M2 ;
			RECT	0 163.735 0.25 163.835 ;
			LAYER	M3 ;
			RECT	0 163.735 0.25 163.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[56]

	PIN QA[57]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 166.615 0.25 166.715 ;
			LAYER	M2 ;
			RECT	0 166.615 0.25 166.715 ;
			LAYER	M3 ;
			RECT	0 166.615 0.25 166.715 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[57]

	PIN QA[58]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 169.495 0.25 169.595 ;
			LAYER	M2 ;
			RECT	0 169.495 0.25 169.595 ;
			LAYER	M3 ;
			RECT	0 169.495 0.25 169.595 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[58]

	PIN QA[59]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 172.375 0.25 172.475 ;
			LAYER	M2 ;
			RECT	0 172.375 0.25 172.475 ;
			LAYER	M3 ;
			RECT	0 172.375 0.25 172.475 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[59]

	PIN QA[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.855 0.25 16.955 ;
			LAYER	M2 ;
			RECT	0 16.855 0.25 16.955 ;
			LAYER	M3 ;
			RECT	0 16.855 0.25 16.955 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[5]

	PIN QA[60]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 175.255 0.25 175.355 ;
			LAYER	M2 ;
			RECT	0 175.255 0.25 175.355 ;
			LAYER	M3 ;
			RECT	0 175.255 0.25 175.355 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[60]

	PIN QA[61]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 178.135 0.25 178.235 ;
			LAYER	M2 ;
			RECT	0 178.135 0.25 178.235 ;
			LAYER	M3 ;
			RECT	0 178.135 0.25 178.235 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[61]

	PIN QA[62]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 181.015 0.25 181.115 ;
			LAYER	M2 ;
			RECT	0 181.015 0.25 181.115 ;
			LAYER	M3 ;
			RECT	0 181.015 0.25 181.115 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[62]

	PIN QA[63]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 183.895 0.25 183.995 ;
			LAYER	M2 ;
			RECT	0 183.895 0.25 183.995 ;
			LAYER	M3 ;
			RECT	0 183.895 0.25 183.995 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[63]

	PIN QA[64]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 230.865 0.25 230.965 ;
			LAYER	M2 ;
			RECT	0 230.865 0.25 230.965 ;
			LAYER	M3 ;
			RECT	0 230.865 0.25 230.965 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[64]

	PIN QA[65]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 233.745 0.25 233.845 ;
			LAYER	M2 ;
			RECT	0 233.745 0.25 233.845 ;
			LAYER	M3 ;
			RECT	0 233.745 0.25 233.845 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[65]

	PIN QA[66]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 236.625 0.25 236.725 ;
			LAYER	M2 ;
			RECT	0 236.625 0.25 236.725 ;
			LAYER	M3 ;
			RECT	0 236.625 0.25 236.725 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[66]

	PIN QA[67]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 239.505 0.25 239.605 ;
			LAYER	M2 ;
			RECT	0 239.505 0.25 239.605 ;
			LAYER	M3 ;
			RECT	0 239.505 0.25 239.605 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[67]

	PIN QA[68]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 242.385 0.25 242.485 ;
			LAYER	M2 ;
			RECT	0 242.385 0.25 242.485 ;
			LAYER	M3 ;
			RECT	0 242.385 0.25 242.485 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[68]

	PIN QA[69]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 245.265 0.25 245.365 ;
			LAYER	M2 ;
			RECT	0 245.265 0.25 245.365 ;
			LAYER	M3 ;
			RECT	0 245.265 0.25 245.365 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[69]

	PIN QA[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.735 0.25 19.835 ;
			LAYER	M2 ;
			RECT	0 19.735 0.25 19.835 ;
			LAYER	M3 ;
			RECT	0 19.735 0.25 19.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[6]

	PIN QA[70]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 248.145 0.25 248.245 ;
			LAYER	M2 ;
			RECT	0 248.145 0.25 248.245 ;
			LAYER	M3 ;
			RECT	0 248.145 0.25 248.245 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[70]

	PIN QA[71]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 251.025 0.25 251.125 ;
			LAYER	M2 ;
			RECT	0 251.025 0.25 251.125 ;
			LAYER	M3 ;
			RECT	0 251.025 0.25 251.125 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[71]

	PIN QA[72]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 253.905 0.25 254.005 ;
			LAYER	M2 ;
			RECT	0 253.905 0.25 254.005 ;
			LAYER	M3 ;
			RECT	0 253.905 0.25 254.005 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[72]

	PIN QA[73]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 256.785 0.25 256.885 ;
			LAYER	M2 ;
			RECT	0 256.785 0.25 256.885 ;
			LAYER	M3 ;
			RECT	0 256.785 0.25 256.885 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[73]

	PIN QA[74]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 259.665 0.25 259.765 ;
			LAYER	M2 ;
			RECT	0 259.665 0.25 259.765 ;
			LAYER	M3 ;
			RECT	0 259.665 0.25 259.765 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[74]

	PIN QA[75]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 262.545 0.25 262.645 ;
			LAYER	M2 ;
			RECT	0 262.545 0.25 262.645 ;
			LAYER	M3 ;
			RECT	0 262.545 0.25 262.645 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[75]

	PIN QA[76]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 265.425 0.25 265.525 ;
			LAYER	M2 ;
			RECT	0 265.425 0.25 265.525 ;
			LAYER	M3 ;
			RECT	0 265.425 0.25 265.525 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[76]

	PIN QA[77]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 268.305 0.25 268.405 ;
			LAYER	M2 ;
			RECT	0 268.305 0.25 268.405 ;
			LAYER	M3 ;
			RECT	0 268.305 0.25 268.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[77]

	PIN QA[78]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 271.185 0.25 271.285 ;
			LAYER	M2 ;
			RECT	0 271.185 0.25 271.285 ;
			LAYER	M3 ;
			RECT	0 271.185 0.25 271.285 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[78]

	PIN QA[79]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 274.065 0.25 274.165 ;
			LAYER	M2 ;
			RECT	0 274.065 0.25 274.165 ;
			LAYER	M3 ;
			RECT	0 274.065 0.25 274.165 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[79]

	PIN QA[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.615 0.25 22.715 ;
			LAYER	M2 ;
			RECT	0 22.615 0.25 22.715 ;
			LAYER	M3 ;
			RECT	0 22.615 0.25 22.715 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[7]

	PIN QA[80]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 276.945 0.25 277.045 ;
			LAYER	M2 ;
			RECT	0 276.945 0.25 277.045 ;
			LAYER	M3 ;
			RECT	0 276.945 0.25 277.045 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[80]

	PIN QA[81]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 279.825 0.25 279.925 ;
			LAYER	M2 ;
			RECT	0 279.825 0.25 279.925 ;
			LAYER	M3 ;
			RECT	0 279.825 0.25 279.925 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[81]

	PIN QA[82]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 282.705 0.25 282.805 ;
			LAYER	M2 ;
			RECT	0 282.705 0.25 282.805 ;
			LAYER	M3 ;
			RECT	0 282.705 0.25 282.805 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[82]

	PIN QA[83]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 285.585 0.25 285.685 ;
			LAYER	M2 ;
			RECT	0 285.585 0.25 285.685 ;
			LAYER	M3 ;
			RECT	0 285.585 0.25 285.685 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[83]

	PIN QA[84]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 288.465 0.25 288.565 ;
			LAYER	M2 ;
			RECT	0 288.465 0.25 288.565 ;
			LAYER	M3 ;
			RECT	0 288.465 0.25 288.565 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[84]

	PIN QA[85]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 291.345 0.25 291.445 ;
			LAYER	M2 ;
			RECT	0 291.345 0.25 291.445 ;
			LAYER	M3 ;
			RECT	0 291.345 0.25 291.445 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[85]

	PIN QA[86]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 294.225 0.25 294.325 ;
			LAYER	M2 ;
			RECT	0 294.225 0.25 294.325 ;
			LAYER	M3 ;
			RECT	0 294.225 0.25 294.325 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[86]

	PIN QA[87]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 297.105 0.25 297.205 ;
			LAYER	M2 ;
			RECT	0 297.105 0.25 297.205 ;
			LAYER	M3 ;
			RECT	0 297.105 0.25 297.205 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[87]

	PIN QA[88]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 299.985 0.25 300.085 ;
			LAYER	M2 ;
			RECT	0 299.985 0.25 300.085 ;
			LAYER	M3 ;
			RECT	0 299.985 0.25 300.085 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[88]

	PIN QA[89]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 302.865 0.25 302.965 ;
			LAYER	M2 ;
			RECT	0 302.865 0.25 302.965 ;
			LAYER	M3 ;
			RECT	0 302.865 0.25 302.965 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[89]

	PIN QA[8]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.495 0.25 25.595 ;
			LAYER	M2 ;
			RECT	0 25.495 0.25 25.595 ;
			LAYER	M3 ;
			RECT	0 25.495 0.25 25.595 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[8]

	PIN QA[90]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 305.745 0.25 305.845 ;
			LAYER	M2 ;
			RECT	0 305.745 0.25 305.845 ;
			LAYER	M3 ;
			RECT	0 305.745 0.25 305.845 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[90]

	PIN QA[91]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 308.625 0.25 308.725 ;
			LAYER	M2 ;
			RECT	0 308.625 0.25 308.725 ;
			LAYER	M3 ;
			RECT	0 308.625 0.25 308.725 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[91]

	PIN QA[92]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 311.505 0.25 311.605 ;
			LAYER	M2 ;
			RECT	0 311.505 0.25 311.605 ;
			LAYER	M3 ;
			RECT	0 311.505 0.25 311.605 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[92]

	PIN QA[93]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 314.385 0.25 314.485 ;
			LAYER	M2 ;
			RECT	0 314.385 0.25 314.485 ;
			LAYER	M3 ;
			RECT	0 314.385 0.25 314.485 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[93]

	PIN QA[94]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 317.265 0.25 317.365 ;
			LAYER	M2 ;
			RECT	0 317.265 0.25 317.365 ;
			LAYER	M3 ;
			RECT	0 317.265 0.25 317.365 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[94]

	PIN QA[95]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 320.145 0.25 320.245 ;
			LAYER	M2 ;
			RECT	0 320.145 0.25 320.245 ;
			LAYER	M3 ;
			RECT	0 320.145 0.25 320.245 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[95]

	PIN QA[96]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 323.025 0.25 323.125 ;
			LAYER	M2 ;
			RECT	0 323.025 0.25 323.125 ;
			LAYER	M3 ;
			RECT	0 323.025 0.25 323.125 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[96]

	PIN QA[97]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 325.905 0.25 326.005 ;
			LAYER	M2 ;
			RECT	0 325.905 0.25 326.005 ;
			LAYER	M3 ;
			RECT	0 325.905 0.25 326.005 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[97]

	PIN QA[98]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 328.785 0.25 328.885 ;
			LAYER	M2 ;
			RECT	0 328.785 0.25 328.885 ;
			LAYER	M3 ;
			RECT	0 328.785 0.25 328.885 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[98]

	PIN QA[99]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 331.665 0.25 331.765 ;
			LAYER	M2 ;
			RECT	0 331.665 0.25 331.765 ;
			LAYER	M3 ;
			RECT	0 331.665 0.25 331.765 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[99]

	PIN QA[9]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 28.375 0.25 28.475 ;
			LAYER	M2 ;
			RECT	0 28.375 0.25 28.475 ;
			LAYER	M3 ;
			RECT	0 28.375 0.25 28.475 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[9]

	PIN RET1N
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 188.11 0.25 188.21 ;
			LAYER	M2 ;
			RECT	0 188.11 0.25 188.21 ;
			LAYER	M3 ;
			RECT	0 188.11 0.25 188.21 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END RET1N

	PIN SEA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 205.9 0.25 206 ;
			LAYER	M2 ;
			RECT	0 205.9 0.25 206 ;
			LAYER	M3 ;
			RECT	0 205.9 0.25 206 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SEA

	PIN SEB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 208.735 0.25 208.835 ;
			LAYER	M2 ;
			RECT	0 208.735 0.25 208.835 ;
			LAYER	M3 ;
			RECT	0 208.735 0.25 208.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SEB

	PIN SIA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 206.1 0.25 206.2 ;
			LAYER	M2 ;
			RECT	0 206.1 0.25 206.2 ;
			LAYER	M3 ;
			RECT	0 206.1 0.25 206.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIA[0]

	PIN SIA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 207.07 0.25 207.17 ;
			LAYER	M2 ;
			RECT	0 207.07 0.25 207.17 ;
			LAYER	M3 ;
			RECT	0 207.07 0.25 207.17 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIA[1]

	PIN SIB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 202.675 0.25 202.775 ;
			LAYER	M2 ;
			RECT	0 202.675 0.25 202.775 ;
			LAYER	M3 ;
			RECT	0 202.675 0.25 202.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIB[0]

	PIN SIB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 220.325 0.25 220.425 ;
			LAYER	M2 ;
			RECT	0 220.325 0.25 220.425 ;
			LAYER	M3 ;
			RECT	0 220.325 0.25 220.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIB[1]

	PIN SOA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 0.36 0.25 0.46 ;
			LAYER	M2 ;
			RECT	0 0.36 0.25 0.46 ;
			LAYER	M3 ;
			RECT	0 0.36 0.25 0.46 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOA[0]

	PIN SOA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 414.4 0.25 414.5 ;
			LAYER	M2 ;
			RECT	0 414.4 0.25 414.5 ;
			LAYER	M3 ;
			RECT	0 414.4 0.25 414.5 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOA[1]

	PIN SOB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 0.09 0.25 0.19 ;
			LAYER	M2 ;
			RECT	0 0.09 0.25 0.19 ;
			LAYER	M3 ;
			RECT	0 0.09 0.25 0.19 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOB[0]

	PIN SOB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 414.67 0.25 414.77 ;
			LAYER	M2 ;
			RECT	0 414.67 0.25 414.77 ;
			LAYER	M3 ;
			RECT	0 414.67 0.25 414.77 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOB[1]

	PIN TAA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 190.755 0.25 190.855 ;
			LAYER	M2 ;
			RECT	0 190.755 0.25 190.855 ;
			LAYER	M3 ;
			RECT	0 190.755 0.25 190.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[0]

	PIN TAA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 193.785 0.25 193.885 ;
			LAYER	M2 ;
			RECT	0 193.785 0.25 193.885 ;
			LAYER	M3 ;
			RECT	0 193.785 0.25 193.885 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[1]

	PIN TAA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 196.845 0.25 196.945 ;
			LAYER	M2 ;
			RECT	0 196.845 0.25 196.945 ;
			LAYER	M3 ;
			RECT	0 196.845 0.25 196.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[2]

	PIN TAA[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 199.36 0.25 199.46 ;
			LAYER	M2 ;
			RECT	0 199.36 0.25 199.46 ;
			LAYER	M3 ;
			RECT	0 199.36 0.25 199.46 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[3]

	PIN TAA[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 202.39 0.25 202.49 ;
			LAYER	M2 ;
			RECT	0 202.39 0.25 202.49 ;
			LAYER	M3 ;
			RECT	0 202.39 0.25 202.49 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[4]

	PIN TAB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 224.67 0.25 224.77 ;
			LAYER	M2 ;
			RECT	0 224.67 0.25 224.77 ;
			LAYER	M3 ;
			RECT	0 224.67 0.25 224.77 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[0]

	PIN TAB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 221.64 0.25 221.74 ;
			LAYER	M2 ;
			RECT	0 221.64 0.25 221.74 ;
			LAYER	M3 ;
			RECT	0 221.64 0.25 221.74 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[1]

	PIN TAB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 218.58 0.25 218.68 ;
			LAYER	M2 ;
			RECT	0 218.58 0.25 218.68 ;
			LAYER	M3 ;
			RECT	0 218.58 0.25 218.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[2]

	PIN TAB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 216.095 0.25 216.195 ;
			LAYER	M2 ;
			RECT	0 216.095 0.25 216.195 ;
			LAYER	M3 ;
			RECT	0 216.095 0.25 216.195 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[3]

	PIN TAB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 213.06 0.25 213.16 ;
			LAYER	M2 ;
			RECT	0 213.06 0.25 213.16 ;
			LAYER	M3 ;
			RECT	0 213.06 0.25 213.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[4]

	PIN TCENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 188.31 0.25 188.41 ;
			LAYER	M2 ;
			RECT	0 188.31 0.25 188.41 ;
			LAYER	M3 ;
			RECT	0 188.31 0.25 188.41 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TCENA

	PIN TCENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 228.31 0.25 228.41 ;
			LAYER	M2 ;
			RECT	0 228.31 0.25 228.41 ;
			LAYER	M3 ;
			RECT	0 228.31 0.25 228.41 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TCENB

	PIN TDB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 1.465 0.25 1.565 ;
			LAYER	M2 ;
			RECT	0 1.465 0.25 1.565 ;
			LAYER	M3 ;
			RECT	0 1.465 0.25 1.565 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[0]

	PIN TDB[100]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 335.535 0.25 335.635 ;
			LAYER	M2 ;
			RECT	0 335.535 0.25 335.635 ;
			LAYER	M3 ;
			RECT	0 335.535 0.25 335.635 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[100]

	PIN TDB[101]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 338.415 0.25 338.515 ;
			LAYER	M2 ;
			RECT	0 338.415 0.25 338.515 ;
			LAYER	M3 ;
			RECT	0 338.415 0.25 338.515 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[101]

	PIN TDB[102]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 341.295 0.25 341.395 ;
			LAYER	M2 ;
			RECT	0 341.295 0.25 341.395 ;
			LAYER	M3 ;
			RECT	0 341.295 0.25 341.395 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[102]

	PIN TDB[103]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 344.175 0.25 344.275 ;
			LAYER	M2 ;
			RECT	0 344.175 0.25 344.275 ;
			LAYER	M3 ;
			RECT	0 344.175 0.25 344.275 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[103]

	PIN TDB[104]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 347.055 0.25 347.155 ;
			LAYER	M2 ;
			RECT	0 347.055 0.25 347.155 ;
			LAYER	M3 ;
			RECT	0 347.055 0.25 347.155 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[104]

	PIN TDB[105]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 349.935 0.25 350.035 ;
			LAYER	M2 ;
			RECT	0 349.935 0.25 350.035 ;
			LAYER	M3 ;
			RECT	0 349.935 0.25 350.035 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[105]

	PIN TDB[106]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 352.815 0.25 352.915 ;
			LAYER	M2 ;
			RECT	0 352.815 0.25 352.915 ;
			LAYER	M3 ;
			RECT	0 352.815 0.25 352.915 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[106]

	PIN TDB[107]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 355.695 0.25 355.795 ;
			LAYER	M2 ;
			RECT	0 355.695 0.25 355.795 ;
			LAYER	M3 ;
			RECT	0 355.695 0.25 355.795 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[107]

	PIN TDB[108]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 358.575 0.25 358.675 ;
			LAYER	M2 ;
			RECT	0 358.575 0.25 358.675 ;
			LAYER	M3 ;
			RECT	0 358.575 0.25 358.675 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[108]

	PIN TDB[109]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 361.455 0.25 361.555 ;
			LAYER	M2 ;
			RECT	0 361.455 0.25 361.555 ;
			LAYER	M3 ;
			RECT	0 361.455 0.25 361.555 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[109]

	PIN TDB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.265 0.25 30.365 ;
			LAYER	M2 ;
			RECT	0 30.265 0.25 30.365 ;
			LAYER	M3 ;
			RECT	0 30.265 0.25 30.365 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[10]

	PIN TDB[110]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 364.335 0.25 364.435 ;
			LAYER	M2 ;
			RECT	0 364.335 0.25 364.435 ;
			LAYER	M3 ;
			RECT	0 364.335 0.25 364.435 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[110]

	PIN TDB[111]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 367.215 0.25 367.315 ;
			LAYER	M2 ;
			RECT	0 367.215 0.25 367.315 ;
			LAYER	M3 ;
			RECT	0 367.215 0.25 367.315 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[111]

	PIN TDB[112]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 370.095 0.25 370.195 ;
			LAYER	M2 ;
			RECT	0 370.095 0.25 370.195 ;
			LAYER	M3 ;
			RECT	0 370.095 0.25 370.195 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[112]

	PIN TDB[113]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 372.975 0.25 373.075 ;
			LAYER	M2 ;
			RECT	0 372.975 0.25 373.075 ;
			LAYER	M3 ;
			RECT	0 372.975 0.25 373.075 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[113]

	PIN TDB[114]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 375.855 0.25 375.955 ;
			LAYER	M2 ;
			RECT	0 375.855 0.25 375.955 ;
			LAYER	M3 ;
			RECT	0 375.855 0.25 375.955 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[114]

	PIN TDB[115]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 378.735 0.25 378.835 ;
			LAYER	M2 ;
			RECT	0 378.735 0.25 378.835 ;
			LAYER	M3 ;
			RECT	0 378.735 0.25 378.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[115]

	PIN TDB[116]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 381.615 0.25 381.715 ;
			LAYER	M2 ;
			RECT	0 381.615 0.25 381.715 ;
			LAYER	M3 ;
			RECT	0 381.615 0.25 381.715 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[116]

	PIN TDB[117]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 384.495 0.25 384.595 ;
			LAYER	M2 ;
			RECT	0 384.495 0.25 384.595 ;
			LAYER	M3 ;
			RECT	0 384.495 0.25 384.595 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[117]

	PIN TDB[118]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 387.375 0.25 387.475 ;
			LAYER	M2 ;
			RECT	0 387.375 0.25 387.475 ;
			LAYER	M3 ;
			RECT	0 387.375 0.25 387.475 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[118]

	PIN TDB[119]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 390.255 0.25 390.355 ;
			LAYER	M2 ;
			RECT	0 390.255 0.25 390.355 ;
			LAYER	M3 ;
			RECT	0 390.255 0.25 390.355 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[119]

	PIN TDB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.145 0.25 33.245 ;
			LAYER	M2 ;
			RECT	0 33.145 0.25 33.245 ;
			LAYER	M3 ;
			RECT	0 33.145 0.25 33.245 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[11]

	PIN TDB[120]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 393.135 0.25 393.235 ;
			LAYER	M2 ;
			RECT	0 393.135 0.25 393.235 ;
			LAYER	M3 ;
			RECT	0 393.135 0.25 393.235 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[120]

	PIN TDB[121]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 396.015 0.25 396.115 ;
			LAYER	M2 ;
			RECT	0 396.015 0.25 396.115 ;
			LAYER	M3 ;
			RECT	0 396.015 0.25 396.115 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[121]

	PIN TDB[122]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 398.895 0.25 398.995 ;
			LAYER	M2 ;
			RECT	0 398.895 0.25 398.995 ;
			LAYER	M3 ;
			RECT	0 398.895 0.25 398.995 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[122]

	PIN TDB[123]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 401.775 0.25 401.875 ;
			LAYER	M2 ;
			RECT	0 401.775 0.25 401.875 ;
			LAYER	M3 ;
			RECT	0 401.775 0.25 401.875 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[123]

	PIN TDB[124]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 404.655 0.25 404.755 ;
			LAYER	M2 ;
			RECT	0 404.655 0.25 404.755 ;
			LAYER	M3 ;
			RECT	0 404.655 0.25 404.755 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[124]

	PIN TDB[125]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 407.535 0.25 407.635 ;
			LAYER	M2 ;
			RECT	0 407.535 0.25 407.635 ;
			LAYER	M3 ;
			RECT	0 407.535 0.25 407.635 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[125]

	PIN TDB[126]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 410.415 0.25 410.515 ;
			LAYER	M2 ;
			RECT	0 410.415 0.25 410.515 ;
			LAYER	M3 ;
			RECT	0 410.415 0.25 410.515 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[126]

	PIN TDB[127]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 413.295 0.25 413.395 ;
			LAYER	M2 ;
			RECT	0 413.295 0.25 413.395 ;
			LAYER	M3 ;
			RECT	0 413.295 0.25 413.395 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[127]

	PIN TDB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.025 0.25 36.125 ;
			LAYER	M2 ;
			RECT	0 36.025 0.25 36.125 ;
			LAYER	M3 ;
			RECT	0 36.025 0.25 36.125 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[12]

	PIN TDB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 38.905 0.25 39.005 ;
			LAYER	M2 ;
			RECT	0 38.905 0.25 39.005 ;
			LAYER	M3 ;
			RECT	0 38.905 0.25 39.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[13]

	PIN TDB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 41.785 0.25 41.885 ;
			LAYER	M2 ;
			RECT	0 41.785 0.25 41.885 ;
			LAYER	M3 ;
			RECT	0 41.785 0.25 41.885 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[14]

	PIN TDB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 44.665 0.25 44.765 ;
			LAYER	M2 ;
			RECT	0 44.665 0.25 44.765 ;
			LAYER	M3 ;
			RECT	0 44.665 0.25 44.765 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[15]

	PIN TDB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.545 0.25 47.645 ;
			LAYER	M2 ;
			RECT	0 47.545 0.25 47.645 ;
			LAYER	M3 ;
			RECT	0 47.545 0.25 47.645 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[16]

	PIN TDB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 50.425 0.25 50.525 ;
			LAYER	M2 ;
			RECT	0 50.425 0.25 50.525 ;
			LAYER	M3 ;
			RECT	0 50.425 0.25 50.525 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[17]

	PIN TDB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 53.305 0.25 53.405 ;
			LAYER	M2 ;
			RECT	0 53.305 0.25 53.405 ;
			LAYER	M3 ;
			RECT	0 53.305 0.25 53.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[18]

	PIN TDB[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.185 0.25 56.285 ;
			LAYER	M2 ;
			RECT	0 56.185 0.25 56.285 ;
			LAYER	M3 ;
			RECT	0 56.185 0.25 56.285 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[19]

	PIN TDB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 4.345 0.25 4.445 ;
			LAYER	M2 ;
			RECT	0 4.345 0.25 4.445 ;
			LAYER	M3 ;
			RECT	0 4.345 0.25 4.445 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[1]

	PIN TDB[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.065 0.25 59.165 ;
			LAYER	M2 ;
			RECT	0 59.065 0.25 59.165 ;
			LAYER	M3 ;
			RECT	0 59.065 0.25 59.165 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[20]

	PIN TDB[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 61.945 0.25 62.045 ;
			LAYER	M2 ;
			RECT	0 61.945 0.25 62.045 ;
			LAYER	M3 ;
			RECT	0 61.945 0.25 62.045 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[21]

	PIN TDB[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 64.825 0.25 64.925 ;
			LAYER	M2 ;
			RECT	0 64.825 0.25 64.925 ;
			LAYER	M3 ;
			RECT	0 64.825 0.25 64.925 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[22]

	PIN TDB[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 67.705 0.25 67.805 ;
			LAYER	M2 ;
			RECT	0 67.705 0.25 67.805 ;
			LAYER	M3 ;
			RECT	0 67.705 0.25 67.805 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[23]

	PIN TDB[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 70.585 0.25 70.685 ;
			LAYER	M2 ;
			RECT	0 70.585 0.25 70.685 ;
			LAYER	M3 ;
			RECT	0 70.585 0.25 70.685 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[24]

	PIN TDB[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 73.465 0.25 73.565 ;
			LAYER	M2 ;
			RECT	0 73.465 0.25 73.565 ;
			LAYER	M3 ;
			RECT	0 73.465 0.25 73.565 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[25]

	PIN TDB[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 76.345 0.25 76.445 ;
			LAYER	M2 ;
			RECT	0 76.345 0.25 76.445 ;
			LAYER	M3 ;
			RECT	0 76.345 0.25 76.445 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[26]

	PIN TDB[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.225 0.25 79.325 ;
			LAYER	M2 ;
			RECT	0 79.225 0.25 79.325 ;
			LAYER	M3 ;
			RECT	0 79.225 0.25 79.325 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[27]

	PIN TDB[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.105 0.25 82.205 ;
			LAYER	M2 ;
			RECT	0 82.105 0.25 82.205 ;
			LAYER	M3 ;
			RECT	0 82.105 0.25 82.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[28]

	PIN TDB[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 84.985 0.25 85.085 ;
			LAYER	M2 ;
			RECT	0 84.985 0.25 85.085 ;
			LAYER	M3 ;
			RECT	0 84.985 0.25 85.085 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[29]

	PIN TDB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.225 0.25 7.325 ;
			LAYER	M2 ;
			RECT	0 7.225 0.25 7.325 ;
			LAYER	M3 ;
			RECT	0 7.225 0.25 7.325 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[2]

	PIN TDB[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 87.865 0.25 87.965 ;
			LAYER	M2 ;
			RECT	0 87.865 0.25 87.965 ;
			LAYER	M3 ;
			RECT	0 87.865 0.25 87.965 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[30]

	PIN TDB[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 90.745 0.25 90.845 ;
			LAYER	M2 ;
			RECT	0 90.745 0.25 90.845 ;
			LAYER	M3 ;
			RECT	0 90.745 0.25 90.845 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[31]

	PIN TDB[32]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 93.625 0.25 93.725 ;
			LAYER	M2 ;
			RECT	0 93.625 0.25 93.725 ;
			LAYER	M3 ;
			RECT	0 93.625 0.25 93.725 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[32]

	PIN TDB[33]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 96.505 0.25 96.605 ;
			LAYER	M2 ;
			RECT	0 96.505 0.25 96.605 ;
			LAYER	M3 ;
			RECT	0 96.505 0.25 96.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[33]

	PIN TDB[34]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 99.385 0.25 99.485 ;
			LAYER	M2 ;
			RECT	0 99.385 0.25 99.485 ;
			LAYER	M3 ;
			RECT	0 99.385 0.25 99.485 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[34]

	PIN TDB[35]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 102.265 0.25 102.365 ;
			LAYER	M2 ;
			RECT	0 102.265 0.25 102.365 ;
			LAYER	M3 ;
			RECT	0 102.265 0.25 102.365 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[35]

	PIN TDB[36]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 105.145 0.25 105.245 ;
			LAYER	M2 ;
			RECT	0 105.145 0.25 105.245 ;
			LAYER	M3 ;
			RECT	0 105.145 0.25 105.245 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[36]

	PIN TDB[37]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 108.025 0.25 108.125 ;
			LAYER	M2 ;
			RECT	0 108.025 0.25 108.125 ;
			LAYER	M3 ;
			RECT	0 108.025 0.25 108.125 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[37]

	PIN TDB[38]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 110.905 0.25 111.005 ;
			LAYER	M2 ;
			RECT	0 110.905 0.25 111.005 ;
			LAYER	M3 ;
			RECT	0 110.905 0.25 111.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[38]

	PIN TDB[39]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 113.785 0.25 113.885 ;
			LAYER	M2 ;
			RECT	0 113.785 0.25 113.885 ;
			LAYER	M3 ;
			RECT	0 113.785 0.25 113.885 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[39]

	PIN TDB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.105 0.25 10.205 ;
			LAYER	M2 ;
			RECT	0 10.105 0.25 10.205 ;
			LAYER	M3 ;
			RECT	0 10.105 0.25 10.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[3]

	PIN TDB[40]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 116.665 0.25 116.765 ;
			LAYER	M2 ;
			RECT	0 116.665 0.25 116.765 ;
			LAYER	M3 ;
			RECT	0 116.665 0.25 116.765 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[40]

	PIN TDB[41]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 119.545 0.25 119.645 ;
			LAYER	M2 ;
			RECT	0 119.545 0.25 119.645 ;
			LAYER	M3 ;
			RECT	0 119.545 0.25 119.645 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[41]

	PIN TDB[42]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 122.425 0.25 122.525 ;
			LAYER	M2 ;
			RECT	0 122.425 0.25 122.525 ;
			LAYER	M3 ;
			RECT	0 122.425 0.25 122.525 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[42]

	PIN TDB[43]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 125.305 0.25 125.405 ;
			LAYER	M2 ;
			RECT	0 125.305 0.25 125.405 ;
			LAYER	M3 ;
			RECT	0 125.305 0.25 125.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[43]

	PIN TDB[44]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 128.185 0.25 128.285 ;
			LAYER	M2 ;
			RECT	0 128.185 0.25 128.285 ;
			LAYER	M3 ;
			RECT	0 128.185 0.25 128.285 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[44]

	PIN TDB[45]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 131.065 0.25 131.165 ;
			LAYER	M2 ;
			RECT	0 131.065 0.25 131.165 ;
			LAYER	M3 ;
			RECT	0 131.065 0.25 131.165 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[45]

	PIN TDB[46]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 133.945 0.25 134.045 ;
			LAYER	M2 ;
			RECT	0 133.945 0.25 134.045 ;
			LAYER	M3 ;
			RECT	0 133.945 0.25 134.045 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[46]

	PIN TDB[47]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 136.825 0.25 136.925 ;
			LAYER	M2 ;
			RECT	0 136.825 0.25 136.925 ;
			LAYER	M3 ;
			RECT	0 136.825 0.25 136.925 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[47]

	PIN TDB[48]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 139.705 0.25 139.805 ;
			LAYER	M2 ;
			RECT	0 139.705 0.25 139.805 ;
			LAYER	M3 ;
			RECT	0 139.705 0.25 139.805 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[48]

	PIN TDB[49]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 142.585 0.25 142.685 ;
			LAYER	M2 ;
			RECT	0 142.585 0.25 142.685 ;
			LAYER	M3 ;
			RECT	0 142.585 0.25 142.685 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[49]

	PIN TDB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 12.985 0.25 13.085 ;
			LAYER	M2 ;
			RECT	0 12.985 0.25 13.085 ;
			LAYER	M3 ;
			RECT	0 12.985 0.25 13.085 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[4]

	PIN TDB[50]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 145.465 0.25 145.565 ;
			LAYER	M2 ;
			RECT	0 145.465 0.25 145.565 ;
			LAYER	M3 ;
			RECT	0 145.465 0.25 145.565 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[50]

	PIN TDB[51]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 148.345 0.25 148.445 ;
			LAYER	M2 ;
			RECT	0 148.345 0.25 148.445 ;
			LAYER	M3 ;
			RECT	0 148.345 0.25 148.445 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[51]

	PIN TDB[52]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 151.225 0.25 151.325 ;
			LAYER	M2 ;
			RECT	0 151.225 0.25 151.325 ;
			LAYER	M3 ;
			RECT	0 151.225 0.25 151.325 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[52]

	PIN TDB[53]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 154.105 0.25 154.205 ;
			LAYER	M2 ;
			RECT	0 154.105 0.25 154.205 ;
			LAYER	M3 ;
			RECT	0 154.105 0.25 154.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[53]

	PIN TDB[54]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 156.985 0.25 157.085 ;
			LAYER	M2 ;
			RECT	0 156.985 0.25 157.085 ;
			LAYER	M3 ;
			RECT	0 156.985 0.25 157.085 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[54]

	PIN TDB[55]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 159.865 0.25 159.965 ;
			LAYER	M2 ;
			RECT	0 159.865 0.25 159.965 ;
			LAYER	M3 ;
			RECT	0 159.865 0.25 159.965 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[55]

	PIN TDB[56]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 162.745 0.25 162.845 ;
			LAYER	M2 ;
			RECT	0 162.745 0.25 162.845 ;
			LAYER	M3 ;
			RECT	0 162.745 0.25 162.845 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[56]

	PIN TDB[57]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 165.625 0.25 165.725 ;
			LAYER	M2 ;
			RECT	0 165.625 0.25 165.725 ;
			LAYER	M3 ;
			RECT	0 165.625 0.25 165.725 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[57]

	PIN TDB[58]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 168.505 0.25 168.605 ;
			LAYER	M2 ;
			RECT	0 168.505 0.25 168.605 ;
			LAYER	M3 ;
			RECT	0 168.505 0.25 168.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[58]

	PIN TDB[59]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 171.385 0.25 171.485 ;
			LAYER	M2 ;
			RECT	0 171.385 0.25 171.485 ;
			LAYER	M3 ;
			RECT	0 171.385 0.25 171.485 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[59]

	PIN TDB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 15.865 0.25 15.965 ;
			LAYER	M2 ;
			RECT	0 15.865 0.25 15.965 ;
			LAYER	M3 ;
			RECT	0 15.865 0.25 15.965 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[5]

	PIN TDB[60]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 174.265 0.25 174.365 ;
			LAYER	M2 ;
			RECT	0 174.265 0.25 174.365 ;
			LAYER	M3 ;
			RECT	0 174.265 0.25 174.365 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[60]

	PIN TDB[61]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 177.145 0.25 177.245 ;
			LAYER	M2 ;
			RECT	0 177.145 0.25 177.245 ;
			LAYER	M3 ;
			RECT	0 177.145 0.25 177.245 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[61]

	PIN TDB[62]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 180.025 0.25 180.125 ;
			LAYER	M2 ;
			RECT	0 180.025 0.25 180.125 ;
			LAYER	M3 ;
			RECT	0 180.025 0.25 180.125 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[62]

	PIN TDB[63]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 182.905 0.25 183.005 ;
			LAYER	M2 ;
			RECT	0 182.905 0.25 183.005 ;
			LAYER	M3 ;
			RECT	0 182.905 0.25 183.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[63]

	PIN TDB[64]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 231.855 0.25 231.955 ;
			LAYER	M2 ;
			RECT	0 231.855 0.25 231.955 ;
			LAYER	M3 ;
			RECT	0 231.855 0.25 231.955 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[64]

	PIN TDB[65]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 234.735 0.25 234.835 ;
			LAYER	M2 ;
			RECT	0 234.735 0.25 234.835 ;
			LAYER	M3 ;
			RECT	0 234.735 0.25 234.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[65]

	PIN TDB[66]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 237.615 0.25 237.715 ;
			LAYER	M2 ;
			RECT	0 237.615 0.25 237.715 ;
			LAYER	M3 ;
			RECT	0 237.615 0.25 237.715 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[66]

	PIN TDB[67]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 240.495 0.25 240.595 ;
			LAYER	M2 ;
			RECT	0 240.495 0.25 240.595 ;
			LAYER	M3 ;
			RECT	0 240.495 0.25 240.595 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[67]

	PIN TDB[68]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 243.375 0.25 243.475 ;
			LAYER	M2 ;
			RECT	0 243.375 0.25 243.475 ;
			LAYER	M3 ;
			RECT	0 243.375 0.25 243.475 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[68]

	PIN TDB[69]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 246.255 0.25 246.355 ;
			LAYER	M2 ;
			RECT	0 246.255 0.25 246.355 ;
			LAYER	M3 ;
			RECT	0 246.255 0.25 246.355 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[69]

	PIN TDB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 18.745 0.25 18.845 ;
			LAYER	M2 ;
			RECT	0 18.745 0.25 18.845 ;
			LAYER	M3 ;
			RECT	0 18.745 0.25 18.845 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[6]

	PIN TDB[70]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 249.135 0.25 249.235 ;
			LAYER	M2 ;
			RECT	0 249.135 0.25 249.235 ;
			LAYER	M3 ;
			RECT	0 249.135 0.25 249.235 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[70]

	PIN TDB[71]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 252.015 0.25 252.115 ;
			LAYER	M2 ;
			RECT	0 252.015 0.25 252.115 ;
			LAYER	M3 ;
			RECT	0 252.015 0.25 252.115 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[71]

	PIN TDB[72]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 254.895 0.25 254.995 ;
			LAYER	M2 ;
			RECT	0 254.895 0.25 254.995 ;
			LAYER	M3 ;
			RECT	0 254.895 0.25 254.995 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[72]

	PIN TDB[73]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 257.775 0.25 257.875 ;
			LAYER	M2 ;
			RECT	0 257.775 0.25 257.875 ;
			LAYER	M3 ;
			RECT	0 257.775 0.25 257.875 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[73]

	PIN TDB[74]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 260.655 0.25 260.755 ;
			LAYER	M2 ;
			RECT	0 260.655 0.25 260.755 ;
			LAYER	M3 ;
			RECT	0 260.655 0.25 260.755 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[74]

	PIN TDB[75]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 263.535 0.25 263.635 ;
			LAYER	M2 ;
			RECT	0 263.535 0.25 263.635 ;
			LAYER	M3 ;
			RECT	0 263.535 0.25 263.635 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[75]

	PIN TDB[76]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 266.415 0.25 266.515 ;
			LAYER	M2 ;
			RECT	0 266.415 0.25 266.515 ;
			LAYER	M3 ;
			RECT	0 266.415 0.25 266.515 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[76]

	PIN TDB[77]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 269.295 0.25 269.395 ;
			LAYER	M2 ;
			RECT	0 269.295 0.25 269.395 ;
			LAYER	M3 ;
			RECT	0 269.295 0.25 269.395 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[77]

	PIN TDB[78]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 272.175 0.25 272.275 ;
			LAYER	M2 ;
			RECT	0 272.175 0.25 272.275 ;
			LAYER	M3 ;
			RECT	0 272.175 0.25 272.275 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[78]

	PIN TDB[79]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 275.055 0.25 275.155 ;
			LAYER	M2 ;
			RECT	0 275.055 0.25 275.155 ;
			LAYER	M3 ;
			RECT	0 275.055 0.25 275.155 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[79]

	PIN TDB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 21.625 0.25 21.725 ;
			LAYER	M2 ;
			RECT	0 21.625 0.25 21.725 ;
			LAYER	M3 ;
			RECT	0 21.625 0.25 21.725 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[7]

	PIN TDB[80]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 277.935 0.25 278.035 ;
			LAYER	M2 ;
			RECT	0 277.935 0.25 278.035 ;
			LAYER	M3 ;
			RECT	0 277.935 0.25 278.035 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[80]

	PIN TDB[81]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 280.815 0.25 280.915 ;
			LAYER	M2 ;
			RECT	0 280.815 0.25 280.915 ;
			LAYER	M3 ;
			RECT	0 280.815 0.25 280.915 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[81]

	PIN TDB[82]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 283.695 0.25 283.795 ;
			LAYER	M2 ;
			RECT	0 283.695 0.25 283.795 ;
			LAYER	M3 ;
			RECT	0 283.695 0.25 283.795 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[82]

	PIN TDB[83]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 286.575 0.25 286.675 ;
			LAYER	M2 ;
			RECT	0 286.575 0.25 286.675 ;
			LAYER	M3 ;
			RECT	0 286.575 0.25 286.675 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[83]

	PIN TDB[84]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 289.455 0.25 289.555 ;
			LAYER	M2 ;
			RECT	0 289.455 0.25 289.555 ;
			LAYER	M3 ;
			RECT	0 289.455 0.25 289.555 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[84]

	PIN TDB[85]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 292.335 0.25 292.435 ;
			LAYER	M2 ;
			RECT	0 292.335 0.25 292.435 ;
			LAYER	M3 ;
			RECT	0 292.335 0.25 292.435 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[85]

	PIN TDB[86]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 295.215 0.25 295.315 ;
			LAYER	M2 ;
			RECT	0 295.215 0.25 295.315 ;
			LAYER	M3 ;
			RECT	0 295.215 0.25 295.315 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[86]

	PIN TDB[87]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 298.095 0.25 298.195 ;
			LAYER	M2 ;
			RECT	0 298.095 0.25 298.195 ;
			LAYER	M3 ;
			RECT	0 298.095 0.25 298.195 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[87]

	PIN TDB[88]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 300.975 0.25 301.075 ;
			LAYER	M2 ;
			RECT	0 300.975 0.25 301.075 ;
			LAYER	M3 ;
			RECT	0 300.975 0.25 301.075 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[88]

	PIN TDB[89]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 303.855 0.25 303.955 ;
			LAYER	M2 ;
			RECT	0 303.855 0.25 303.955 ;
			LAYER	M3 ;
			RECT	0 303.855 0.25 303.955 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[89]

	PIN TDB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 24.505 0.25 24.605 ;
			LAYER	M2 ;
			RECT	0 24.505 0.25 24.605 ;
			LAYER	M3 ;
			RECT	0 24.505 0.25 24.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[8]

	PIN TDB[90]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 306.735 0.25 306.835 ;
			LAYER	M2 ;
			RECT	0 306.735 0.25 306.835 ;
			LAYER	M3 ;
			RECT	0 306.735 0.25 306.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[90]

	PIN TDB[91]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 309.615 0.25 309.715 ;
			LAYER	M2 ;
			RECT	0 309.615 0.25 309.715 ;
			LAYER	M3 ;
			RECT	0 309.615 0.25 309.715 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[91]

	PIN TDB[92]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 312.495 0.25 312.595 ;
			LAYER	M2 ;
			RECT	0 312.495 0.25 312.595 ;
			LAYER	M3 ;
			RECT	0 312.495 0.25 312.595 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[92]

	PIN TDB[93]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 315.375 0.25 315.475 ;
			LAYER	M2 ;
			RECT	0 315.375 0.25 315.475 ;
			LAYER	M3 ;
			RECT	0 315.375 0.25 315.475 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[93]

	PIN TDB[94]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 318.255 0.25 318.355 ;
			LAYER	M2 ;
			RECT	0 318.255 0.25 318.355 ;
			LAYER	M3 ;
			RECT	0 318.255 0.25 318.355 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[94]

	PIN TDB[95]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 321.135 0.25 321.235 ;
			LAYER	M2 ;
			RECT	0 321.135 0.25 321.235 ;
			LAYER	M3 ;
			RECT	0 321.135 0.25 321.235 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[95]

	PIN TDB[96]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 324.015 0.25 324.115 ;
			LAYER	M2 ;
			RECT	0 324.015 0.25 324.115 ;
			LAYER	M3 ;
			RECT	0 324.015 0.25 324.115 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[96]

	PIN TDB[97]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 326.895 0.25 326.995 ;
			LAYER	M2 ;
			RECT	0 326.895 0.25 326.995 ;
			LAYER	M3 ;
			RECT	0 326.895 0.25 326.995 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[97]

	PIN TDB[98]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 329.775 0.25 329.875 ;
			LAYER	M2 ;
			RECT	0 329.775 0.25 329.875 ;
			LAYER	M3 ;
			RECT	0 329.775 0.25 329.875 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[98]

	PIN TDB[99]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 332.655 0.25 332.755 ;
			LAYER	M2 ;
			RECT	0 332.655 0.25 332.755 ;
			LAYER	M3 ;
			RECT	0 332.655 0.25 332.755 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[99]

	PIN TDB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 27.385 0.25 27.485 ;
			LAYER	M2 ;
			RECT	0 27.385 0.25 27.485 ;
			LAYER	M3 ;
			RECT	0 27.385 0.25 27.485 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[9]

	PIN TENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 190.45 0.25 190.55 ;
			LAYER	M2 ;
			RECT	0 190.45 0.25 190.55 ;
			LAYER	M3 ;
			RECT	0 190.45 0.25 190.55 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TENA

	PIN TENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 224.925 0.25 225.025 ;
			LAYER	M2 ;
			RECT	0 224.925 0.25 225.025 ;
			LAYER	M3 ;
			RECT	0 224.925 0.25 225.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TENB

	PIN TWENB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 3.26 0.25 3.36 ;
			LAYER	M2 ;
			RECT	0 3.26 0.25 3.36 ;
			LAYER	M3 ;
			RECT	0 3.26 0.25 3.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[0]

	PIN TWENB[100]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 333.74 0.25 333.84 ;
			LAYER	M2 ;
			RECT	0 333.74 0.25 333.84 ;
			LAYER	M3 ;
			RECT	0 333.74 0.25 333.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[100]

	PIN TWENB[101]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 336.62 0.25 336.72 ;
			LAYER	M2 ;
			RECT	0 336.62 0.25 336.72 ;
			LAYER	M3 ;
			RECT	0 336.62 0.25 336.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[101]

	PIN TWENB[102]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 339.5 0.25 339.6 ;
			LAYER	M2 ;
			RECT	0 339.5 0.25 339.6 ;
			LAYER	M3 ;
			RECT	0 339.5 0.25 339.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[102]

	PIN TWENB[103]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 342.38 0.25 342.48 ;
			LAYER	M2 ;
			RECT	0 342.38 0.25 342.48 ;
			LAYER	M3 ;
			RECT	0 342.38 0.25 342.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[103]

	PIN TWENB[104]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 345.26 0.25 345.36 ;
			LAYER	M2 ;
			RECT	0 345.26 0.25 345.36 ;
			LAYER	M3 ;
			RECT	0 345.26 0.25 345.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[104]

	PIN TWENB[105]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 348.14 0.25 348.24 ;
			LAYER	M2 ;
			RECT	0 348.14 0.25 348.24 ;
			LAYER	M3 ;
			RECT	0 348.14 0.25 348.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[105]

	PIN TWENB[106]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 351.02 0.25 351.12 ;
			LAYER	M2 ;
			RECT	0 351.02 0.25 351.12 ;
			LAYER	M3 ;
			RECT	0 351.02 0.25 351.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[106]

	PIN TWENB[107]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 353.9 0.25 354 ;
			LAYER	M2 ;
			RECT	0 353.9 0.25 354 ;
			LAYER	M3 ;
			RECT	0 353.9 0.25 354 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[107]

	PIN TWENB[108]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 356.78 0.25 356.88 ;
			LAYER	M2 ;
			RECT	0 356.78 0.25 356.88 ;
			LAYER	M3 ;
			RECT	0 356.78 0.25 356.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[108]

	PIN TWENB[109]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 359.66 0.25 359.76 ;
			LAYER	M2 ;
			RECT	0 359.66 0.25 359.76 ;
			LAYER	M3 ;
			RECT	0 359.66 0.25 359.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[109]

	PIN TWENB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 32.06 0.25 32.16 ;
			LAYER	M2 ;
			RECT	0 32.06 0.25 32.16 ;
			LAYER	M3 ;
			RECT	0 32.06 0.25 32.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[10]

	PIN TWENB[110]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 362.54 0.25 362.64 ;
			LAYER	M2 ;
			RECT	0 362.54 0.25 362.64 ;
			LAYER	M3 ;
			RECT	0 362.54 0.25 362.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[110]

	PIN TWENB[111]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 365.42 0.25 365.52 ;
			LAYER	M2 ;
			RECT	0 365.42 0.25 365.52 ;
			LAYER	M3 ;
			RECT	0 365.42 0.25 365.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[111]

	PIN TWENB[112]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 368.3 0.25 368.4 ;
			LAYER	M2 ;
			RECT	0 368.3 0.25 368.4 ;
			LAYER	M3 ;
			RECT	0 368.3 0.25 368.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[112]

	PIN TWENB[113]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 371.18 0.25 371.28 ;
			LAYER	M2 ;
			RECT	0 371.18 0.25 371.28 ;
			LAYER	M3 ;
			RECT	0 371.18 0.25 371.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[113]

	PIN TWENB[114]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 374.06 0.25 374.16 ;
			LAYER	M2 ;
			RECT	0 374.06 0.25 374.16 ;
			LAYER	M3 ;
			RECT	0 374.06 0.25 374.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[114]

	PIN TWENB[115]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 376.94 0.25 377.04 ;
			LAYER	M2 ;
			RECT	0 376.94 0.25 377.04 ;
			LAYER	M3 ;
			RECT	0 376.94 0.25 377.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[115]

	PIN TWENB[116]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 379.82 0.25 379.92 ;
			LAYER	M2 ;
			RECT	0 379.82 0.25 379.92 ;
			LAYER	M3 ;
			RECT	0 379.82 0.25 379.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[116]

	PIN TWENB[117]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 382.7 0.25 382.8 ;
			LAYER	M2 ;
			RECT	0 382.7 0.25 382.8 ;
			LAYER	M3 ;
			RECT	0 382.7 0.25 382.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[117]

	PIN TWENB[118]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 385.58 0.25 385.68 ;
			LAYER	M2 ;
			RECT	0 385.58 0.25 385.68 ;
			LAYER	M3 ;
			RECT	0 385.58 0.25 385.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[118]

	PIN TWENB[119]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 388.46 0.25 388.56 ;
			LAYER	M2 ;
			RECT	0 388.46 0.25 388.56 ;
			LAYER	M3 ;
			RECT	0 388.46 0.25 388.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[119]

	PIN TWENB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 34.94 0.25 35.04 ;
			LAYER	M2 ;
			RECT	0 34.94 0.25 35.04 ;
			LAYER	M3 ;
			RECT	0 34.94 0.25 35.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[11]

	PIN TWENB[120]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 391.34 0.25 391.44 ;
			LAYER	M2 ;
			RECT	0 391.34 0.25 391.44 ;
			LAYER	M3 ;
			RECT	0 391.34 0.25 391.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[120]

	PIN TWENB[121]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 394.22 0.25 394.32 ;
			LAYER	M2 ;
			RECT	0 394.22 0.25 394.32 ;
			LAYER	M3 ;
			RECT	0 394.22 0.25 394.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[121]

	PIN TWENB[122]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 397.1 0.25 397.2 ;
			LAYER	M2 ;
			RECT	0 397.1 0.25 397.2 ;
			LAYER	M3 ;
			RECT	0 397.1 0.25 397.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[122]

	PIN TWENB[123]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 399.98 0.25 400.08 ;
			LAYER	M2 ;
			RECT	0 399.98 0.25 400.08 ;
			LAYER	M3 ;
			RECT	0 399.98 0.25 400.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[123]

	PIN TWENB[124]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 402.86 0.25 402.96 ;
			LAYER	M2 ;
			RECT	0 402.86 0.25 402.96 ;
			LAYER	M3 ;
			RECT	0 402.86 0.25 402.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[124]

	PIN TWENB[125]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 405.74 0.25 405.84 ;
			LAYER	M2 ;
			RECT	0 405.74 0.25 405.84 ;
			LAYER	M3 ;
			RECT	0 405.74 0.25 405.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[125]

	PIN TWENB[126]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 408.62 0.25 408.72 ;
			LAYER	M2 ;
			RECT	0 408.62 0.25 408.72 ;
			LAYER	M3 ;
			RECT	0 408.62 0.25 408.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[126]

	PIN TWENB[127]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 411.5 0.25 411.6 ;
			LAYER	M2 ;
			RECT	0 411.5 0.25 411.6 ;
			LAYER	M3 ;
			RECT	0 411.5 0.25 411.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[127]

	PIN TWENB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 37.82 0.25 37.92 ;
			LAYER	M2 ;
			RECT	0 37.82 0.25 37.92 ;
			LAYER	M3 ;
			RECT	0 37.82 0.25 37.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[12]

	PIN TWENB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 40.7 0.25 40.8 ;
			LAYER	M2 ;
			RECT	0 40.7 0.25 40.8 ;
			LAYER	M3 ;
			RECT	0 40.7 0.25 40.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[13]

	PIN TWENB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.58 0.25 43.68 ;
			LAYER	M2 ;
			RECT	0 43.58 0.25 43.68 ;
			LAYER	M3 ;
			RECT	0 43.58 0.25 43.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[14]

	PIN TWENB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 46.46 0.25 46.56 ;
			LAYER	M2 ;
			RECT	0 46.46 0.25 46.56 ;
			LAYER	M3 ;
			RECT	0 46.46 0.25 46.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[15]

	PIN TWENB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 49.34 0.25 49.44 ;
			LAYER	M2 ;
			RECT	0 49.34 0.25 49.44 ;
			LAYER	M3 ;
			RECT	0 49.34 0.25 49.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[16]

	PIN TWENB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 52.22 0.25 52.32 ;
			LAYER	M2 ;
			RECT	0 52.22 0.25 52.32 ;
			LAYER	M3 ;
			RECT	0 52.22 0.25 52.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[17]

	PIN TWENB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 55.1 0.25 55.2 ;
			LAYER	M2 ;
			RECT	0 55.1 0.25 55.2 ;
			LAYER	M3 ;
			RECT	0 55.1 0.25 55.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[18]

	PIN TWENB[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 57.98 0.25 58.08 ;
			LAYER	M2 ;
			RECT	0 57.98 0.25 58.08 ;
			LAYER	M3 ;
			RECT	0 57.98 0.25 58.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[19]

	PIN TWENB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 6.14 0.25 6.24 ;
			LAYER	M2 ;
			RECT	0 6.14 0.25 6.24 ;
			LAYER	M3 ;
			RECT	0 6.14 0.25 6.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[1]

	PIN TWENB[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.86 0.25 60.96 ;
			LAYER	M2 ;
			RECT	0 60.86 0.25 60.96 ;
			LAYER	M3 ;
			RECT	0 60.86 0.25 60.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[20]

	PIN TWENB[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 63.74 0.25 63.84 ;
			LAYER	M2 ;
			RECT	0 63.74 0.25 63.84 ;
			LAYER	M3 ;
			RECT	0 63.74 0.25 63.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[21]

	PIN TWENB[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 66.62 0.25 66.72 ;
			LAYER	M2 ;
			RECT	0 66.62 0.25 66.72 ;
			LAYER	M3 ;
			RECT	0 66.62 0.25 66.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[22]

	PIN TWENB[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 69.5 0.25 69.6 ;
			LAYER	M2 ;
			RECT	0 69.5 0.25 69.6 ;
			LAYER	M3 ;
			RECT	0 69.5 0.25 69.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[23]

	PIN TWENB[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 72.38 0.25 72.48 ;
			LAYER	M2 ;
			RECT	0 72.38 0.25 72.48 ;
			LAYER	M3 ;
			RECT	0 72.38 0.25 72.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[24]

	PIN TWENB[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 75.26 0.25 75.36 ;
			LAYER	M2 ;
			RECT	0 75.26 0.25 75.36 ;
			LAYER	M3 ;
			RECT	0 75.26 0.25 75.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[25]

	PIN TWENB[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 78.14 0.25 78.24 ;
			LAYER	M2 ;
			RECT	0 78.14 0.25 78.24 ;
			LAYER	M3 ;
			RECT	0 78.14 0.25 78.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[26]

	PIN TWENB[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 81.02 0.25 81.12 ;
			LAYER	M2 ;
			RECT	0 81.02 0.25 81.12 ;
			LAYER	M3 ;
			RECT	0 81.02 0.25 81.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[27]

	PIN TWENB[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 83.9 0.25 84 ;
			LAYER	M2 ;
			RECT	0 83.9 0.25 84 ;
			LAYER	M3 ;
			RECT	0 83.9 0.25 84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[28]

	PIN TWENB[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 86.78 0.25 86.88 ;
			LAYER	M2 ;
			RECT	0 86.78 0.25 86.88 ;
			LAYER	M3 ;
			RECT	0 86.78 0.25 86.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[29]

	PIN TWENB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 9.02 0.25 9.12 ;
			LAYER	M2 ;
			RECT	0 9.02 0.25 9.12 ;
			LAYER	M3 ;
			RECT	0 9.02 0.25 9.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[2]

	PIN TWENB[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 89.66 0.25 89.76 ;
			LAYER	M2 ;
			RECT	0 89.66 0.25 89.76 ;
			LAYER	M3 ;
			RECT	0 89.66 0.25 89.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[30]

	PIN TWENB[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 92.54 0.25 92.64 ;
			LAYER	M2 ;
			RECT	0 92.54 0.25 92.64 ;
			LAYER	M3 ;
			RECT	0 92.54 0.25 92.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[31]

	PIN TWENB[32]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 95.42 0.25 95.52 ;
			LAYER	M2 ;
			RECT	0 95.42 0.25 95.52 ;
			LAYER	M3 ;
			RECT	0 95.42 0.25 95.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[32]

	PIN TWENB[33]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 98.3 0.25 98.4 ;
			LAYER	M2 ;
			RECT	0 98.3 0.25 98.4 ;
			LAYER	M3 ;
			RECT	0 98.3 0.25 98.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[33]

	PIN TWENB[34]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 101.18 0.25 101.28 ;
			LAYER	M2 ;
			RECT	0 101.18 0.25 101.28 ;
			LAYER	M3 ;
			RECT	0 101.18 0.25 101.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[34]

	PIN TWENB[35]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 104.06 0.25 104.16 ;
			LAYER	M2 ;
			RECT	0 104.06 0.25 104.16 ;
			LAYER	M3 ;
			RECT	0 104.06 0.25 104.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[35]

	PIN TWENB[36]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 106.94 0.25 107.04 ;
			LAYER	M2 ;
			RECT	0 106.94 0.25 107.04 ;
			LAYER	M3 ;
			RECT	0 106.94 0.25 107.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[36]

	PIN TWENB[37]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 109.82 0.25 109.92 ;
			LAYER	M2 ;
			RECT	0 109.82 0.25 109.92 ;
			LAYER	M3 ;
			RECT	0 109.82 0.25 109.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[37]

	PIN TWENB[38]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 112.7 0.25 112.8 ;
			LAYER	M2 ;
			RECT	0 112.7 0.25 112.8 ;
			LAYER	M3 ;
			RECT	0 112.7 0.25 112.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[38]

	PIN TWENB[39]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 115.58 0.25 115.68 ;
			LAYER	M2 ;
			RECT	0 115.58 0.25 115.68 ;
			LAYER	M3 ;
			RECT	0 115.58 0.25 115.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[39]

	PIN TWENB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 11.9 0.25 12 ;
			LAYER	M2 ;
			RECT	0 11.9 0.25 12 ;
			LAYER	M3 ;
			RECT	0 11.9 0.25 12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[3]

	PIN TWENB[40]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 118.46 0.25 118.56 ;
			LAYER	M2 ;
			RECT	0 118.46 0.25 118.56 ;
			LAYER	M3 ;
			RECT	0 118.46 0.25 118.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[40]

	PIN TWENB[41]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 121.34 0.25 121.44 ;
			LAYER	M2 ;
			RECT	0 121.34 0.25 121.44 ;
			LAYER	M3 ;
			RECT	0 121.34 0.25 121.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[41]

	PIN TWENB[42]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 124.22 0.25 124.32 ;
			LAYER	M2 ;
			RECT	0 124.22 0.25 124.32 ;
			LAYER	M3 ;
			RECT	0 124.22 0.25 124.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[42]

	PIN TWENB[43]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 127.1 0.25 127.2 ;
			LAYER	M2 ;
			RECT	0 127.1 0.25 127.2 ;
			LAYER	M3 ;
			RECT	0 127.1 0.25 127.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[43]

	PIN TWENB[44]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 129.98 0.25 130.08 ;
			LAYER	M2 ;
			RECT	0 129.98 0.25 130.08 ;
			LAYER	M3 ;
			RECT	0 129.98 0.25 130.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[44]

	PIN TWENB[45]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 132.86 0.25 132.96 ;
			LAYER	M2 ;
			RECT	0 132.86 0.25 132.96 ;
			LAYER	M3 ;
			RECT	0 132.86 0.25 132.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[45]

	PIN TWENB[46]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 135.74 0.25 135.84 ;
			LAYER	M2 ;
			RECT	0 135.74 0.25 135.84 ;
			LAYER	M3 ;
			RECT	0 135.74 0.25 135.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[46]

	PIN TWENB[47]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 138.62 0.25 138.72 ;
			LAYER	M2 ;
			RECT	0 138.62 0.25 138.72 ;
			LAYER	M3 ;
			RECT	0 138.62 0.25 138.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[47]

	PIN TWENB[48]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 141.5 0.25 141.6 ;
			LAYER	M2 ;
			RECT	0 141.5 0.25 141.6 ;
			LAYER	M3 ;
			RECT	0 141.5 0.25 141.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[48]

	PIN TWENB[49]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 144.38 0.25 144.48 ;
			LAYER	M2 ;
			RECT	0 144.38 0.25 144.48 ;
			LAYER	M3 ;
			RECT	0 144.38 0.25 144.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[49]

	PIN TWENB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 14.78 0.25 14.88 ;
			LAYER	M2 ;
			RECT	0 14.78 0.25 14.88 ;
			LAYER	M3 ;
			RECT	0 14.78 0.25 14.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[4]

	PIN TWENB[50]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 147.26 0.25 147.36 ;
			LAYER	M2 ;
			RECT	0 147.26 0.25 147.36 ;
			LAYER	M3 ;
			RECT	0 147.26 0.25 147.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[50]

	PIN TWENB[51]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 150.14 0.25 150.24 ;
			LAYER	M2 ;
			RECT	0 150.14 0.25 150.24 ;
			LAYER	M3 ;
			RECT	0 150.14 0.25 150.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[51]

	PIN TWENB[52]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 153.02 0.25 153.12 ;
			LAYER	M2 ;
			RECT	0 153.02 0.25 153.12 ;
			LAYER	M3 ;
			RECT	0 153.02 0.25 153.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[52]

	PIN TWENB[53]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 155.9 0.25 156 ;
			LAYER	M2 ;
			RECT	0 155.9 0.25 156 ;
			LAYER	M3 ;
			RECT	0 155.9 0.25 156 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[53]

	PIN TWENB[54]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 158.78 0.25 158.88 ;
			LAYER	M2 ;
			RECT	0 158.78 0.25 158.88 ;
			LAYER	M3 ;
			RECT	0 158.78 0.25 158.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[54]

	PIN TWENB[55]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 161.66 0.25 161.76 ;
			LAYER	M2 ;
			RECT	0 161.66 0.25 161.76 ;
			LAYER	M3 ;
			RECT	0 161.66 0.25 161.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[55]

	PIN TWENB[56]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 164.54 0.25 164.64 ;
			LAYER	M2 ;
			RECT	0 164.54 0.25 164.64 ;
			LAYER	M3 ;
			RECT	0 164.54 0.25 164.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[56]

	PIN TWENB[57]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 167.42 0.25 167.52 ;
			LAYER	M2 ;
			RECT	0 167.42 0.25 167.52 ;
			LAYER	M3 ;
			RECT	0 167.42 0.25 167.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[57]

	PIN TWENB[58]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 170.3 0.25 170.4 ;
			LAYER	M2 ;
			RECT	0 170.3 0.25 170.4 ;
			LAYER	M3 ;
			RECT	0 170.3 0.25 170.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[58]

	PIN TWENB[59]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 173.18 0.25 173.28 ;
			LAYER	M2 ;
			RECT	0 173.18 0.25 173.28 ;
			LAYER	M3 ;
			RECT	0 173.18 0.25 173.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[59]

	PIN TWENB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 17.66 0.25 17.76 ;
			LAYER	M2 ;
			RECT	0 17.66 0.25 17.76 ;
			LAYER	M3 ;
			RECT	0 17.66 0.25 17.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[5]

	PIN TWENB[60]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 176.06 0.25 176.16 ;
			LAYER	M2 ;
			RECT	0 176.06 0.25 176.16 ;
			LAYER	M3 ;
			RECT	0 176.06 0.25 176.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[60]

	PIN TWENB[61]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 178.94 0.25 179.04 ;
			LAYER	M2 ;
			RECT	0 178.94 0.25 179.04 ;
			LAYER	M3 ;
			RECT	0 178.94 0.25 179.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[61]

	PIN TWENB[62]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 181.82 0.25 181.92 ;
			LAYER	M2 ;
			RECT	0 181.82 0.25 181.92 ;
			LAYER	M3 ;
			RECT	0 181.82 0.25 181.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[62]

	PIN TWENB[63]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 184.7 0.25 184.8 ;
			LAYER	M2 ;
			RECT	0 184.7 0.25 184.8 ;
			LAYER	M3 ;
			RECT	0 184.7 0.25 184.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[63]

	PIN TWENB[64]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 230.06 0.25 230.16 ;
			LAYER	M2 ;
			RECT	0 230.06 0.25 230.16 ;
			LAYER	M3 ;
			RECT	0 230.06 0.25 230.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[64]

	PIN TWENB[65]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 232.94 0.25 233.04 ;
			LAYER	M2 ;
			RECT	0 232.94 0.25 233.04 ;
			LAYER	M3 ;
			RECT	0 232.94 0.25 233.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[65]

	PIN TWENB[66]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 235.82 0.25 235.92 ;
			LAYER	M2 ;
			RECT	0 235.82 0.25 235.92 ;
			LAYER	M3 ;
			RECT	0 235.82 0.25 235.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[66]

	PIN TWENB[67]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 238.7 0.25 238.8 ;
			LAYER	M2 ;
			RECT	0 238.7 0.25 238.8 ;
			LAYER	M3 ;
			RECT	0 238.7 0.25 238.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[67]

	PIN TWENB[68]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 241.58 0.25 241.68 ;
			LAYER	M2 ;
			RECT	0 241.58 0.25 241.68 ;
			LAYER	M3 ;
			RECT	0 241.58 0.25 241.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[68]

	PIN TWENB[69]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 244.46 0.25 244.56 ;
			LAYER	M2 ;
			RECT	0 244.46 0.25 244.56 ;
			LAYER	M3 ;
			RECT	0 244.46 0.25 244.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[69]

	PIN TWENB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 20.54 0.25 20.64 ;
			LAYER	M2 ;
			RECT	0 20.54 0.25 20.64 ;
			LAYER	M3 ;
			RECT	0 20.54 0.25 20.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[6]

	PIN TWENB[70]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 247.34 0.25 247.44 ;
			LAYER	M2 ;
			RECT	0 247.34 0.25 247.44 ;
			LAYER	M3 ;
			RECT	0 247.34 0.25 247.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[70]

	PIN TWENB[71]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 250.22 0.25 250.32 ;
			LAYER	M2 ;
			RECT	0 250.22 0.25 250.32 ;
			LAYER	M3 ;
			RECT	0 250.22 0.25 250.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[71]

	PIN TWENB[72]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 253.1 0.25 253.2 ;
			LAYER	M2 ;
			RECT	0 253.1 0.25 253.2 ;
			LAYER	M3 ;
			RECT	0 253.1 0.25 253.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[72]

	PIN TWENB[73]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 255.98 0.25 256.08 ;
			LAYER	M2 ;
			RECT	0 255.98 0.25 256.08 ;
			LAYER	M3 ;
			RECT	0 255.98 0.25 256.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[73]

	PIN TWENB[74]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 258.86 0.25 258.96 ;
			LAYER	M2 ;
			RECT	0 258.86 0.25 258.96 ;
			LAYER	M3 ;
			RECT	0 258.86 0.25 258.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[74]

	PIN TWENB[75]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 261.74 0.25 261.84 ;
			LAYER	M2 ;
			RECT	0 261.74 0.25 261.84 ;
			LAYER	M3 ;
			RECT	0 261.74 0.25 261.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[75]

	PIN TWENB[76]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 264.62 0.25 264.72 ;
			LAYER	M2 ;
			RECT	0 264.62 0.25 264.72 ;
			LAYER	M3 ;
			RECT	0 264.62 0.25 264.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[76]

	PIN TWENB[77]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 267.5 0.25 267.6 ;
			LAYER	M2 ;
			RECT	0 267.5 0.25 267.6 ;
			LAYER	M3 ;
			RECT	0 267.5 0.25 267.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[77]

	PIN TWENB[78]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 270.38 0.25 270.48 ;
			LAYER	M2 ;
			RECT	0 270.38 0.25 270.48 ;
			LAYER	M3 ;
			RECT	0 270.38 0.25 270.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[78]

	PIN TWENB[79]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 273.26 0.25 273.36 ;
			LAYER	M2 ;
			RECT	0 273.26 0.25 273.36 ;
			LAYER	M3 ;
			RECT	0 273.26 0.25 273.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[79]

	PIN TWENB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 23.42 0.25 23.52 ;
			LAYER	M2 ;
			RECT	0 23.42 0.25 23.52 ;
			LAYER	M3 ;
			RECT	0 23.42 0.25 23.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[7]

	PIN TWENB[80]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 276.14 0.25 276.24 ;
			LAYER	M2 ;
			RECT	0 276.14 0.25 276.24 ;
			LAYER	M3 ;
			RECT	0 276.14 0.25 276.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[80]

	PIN TWENB[81]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 279.02 0.25 279.12 ;
			LAYER	M2 ;
			RECT	0 279.02 0.25 279.12 ;
			LAYER	M3 ;
			RECT	0 279.02 0.25 279.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[81]

	PIN TWENB[82]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 281.9 0.25 282 ;
			LAYER	M2 ;
			RECT	0 281.9 0.25 282 ;
			LAYER	M3 ;
			RECT	0 281.9 0.25 282 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[82]

	PIN TWENB[83]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 284.78 0.25 284.88 ;
			LAYER	M2 ;
			RECT	0 284.78 0.25 284.88 ;
			LAYER	M3 ;
			RECT	0 284.78 0.25 284.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[83]

	PIN TWENB[84]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 287.66 0.25 287.76 ;
			LAYER	M2 ;
			RECT	0 287.66 0.25 287.76 ;
			LAYER	M3 ;
			RECT	0 287.66 0.25 287.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[84]

	PIN TWENB[85]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 290.54 0.25 290.64 ;
			LAYER	M2 ;
			RECT	0 290.54 0.25 290.64 ;
			LAYER	M3 ;
			RECT	0 290.54 0.25 290.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[85]

	PIN TWENB[86]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 293.42 0.25 293.52 ;
			LAYER	M2 ;
			RECT	0 293.42 0.25 293.52 ;
			LAYER	M3 ;
			RECT	0 293.42 0.25 293.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[86]

	PIN TWENB[87]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 296.3 0.25 296.4 ;
			LAYER	M2 ;
			RECT	0 296.3 0.25 296.4 ;
			LAYER	M3 ;
			RECT	0 296.3 0.25 296.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[87]

	PIN TWENB[88]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 299.18 0.25 299.28 ;
			LAYER	M2 ;
			RECT	0 299.18 0.25 299.28 ;
			LAYER	M3 ;
			RECT	0 299.18 0.25 299.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[88]

	PIN TWENB[89]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 302.06 0.25 302.16 ;
			LAYER	M2 ;
			RECT	0 302.06 0.25 302.16 ;
			LAYER	M3 ;
			RECT	0 302.06 0.25 302.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[89]

	PIN TWENB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 26.3 0.25 26.4 ;
			LAYER	M2 ;
			RECT	0 26.3 0.25 26.4 ;
			LAYER	M3 ;
			RECT	0 26.3 0.25 26.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[8]

	PIN TWENB[90]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 304.94 0.25 305.04 ;
			LAYER	M2 ;
			RECT	0 304.94 0.25 305.04 ;
			LAYER	M3 ;
			RECT	0 304.94 0.25 305.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[90]

	PIN TWENB[91]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 307.82 0.25 307.92 ;
			LAYER	M2 ;
			RECT	0 307.82 0.25 307.92 ;
			LAYER	M3 ;
			RECT	0 307.82 0.25 307.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[91]

	PIN TWENB[92]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 310.7 0.25 310.8 ;
			LAYER	M2 ;
			RECT	0 310.7 0.25 310.8 ;
			LAYER	M3 ;
			RECT	0 310.7 0.25 310.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[92]

	PIN TWENB[93]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 313.58 0.25 313.68 ;
			LAYER	M2 ;
			RECT	0 313.58 0.25 313.68 ;
			LAYER	M3 ;
			RECT	0 313.58 0.25 313.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[93]

	PIN TWENB[94]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 316.46 0.25 316.56 ;
			LAYER	M2 ;
			RECT	0 316.46 0.25 316.56 ;
			LAYER	M3 ;
			RECT	0 316.46 0.25 316.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[94]

	PIN TWENB[95]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 319.34 0.25 319.44 ;
			LAYER	M2 ;
			RECT	0 319.34 0.25 319.44 ;
			LAYER	M3 ;
			RECT	0 319.34 0.25 319.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[95]

	PIN TWENB[96]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 322.22 0.25 322.32 ;
			LAYER	M2 ;
			RECT	0 322.22 0.25 322.32 ;
			LAYER	M3 ;
			RECT	0 322.22 0.25 322.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[96]

	PIN TWENB[97]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 325.1 0.25 325.2 ;
			LAYER	M2 ;
			RECT	0 325.1 0.25 325.2 ;
			LAYER	M3 ;
			RECT	0 325.1 0.25 325.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[97]

	PIN TWENB[98]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 327.98 0.25 328.08 ;
			LAYER	M2 ;
			RECT	0 327.98 0.25 328.08 ;
			LAYER	M3 ;
			RECT	0 327.98 0.25 328.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[98]

	PIN TWENB[99]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 330.86 0.25 330.96 ;
			LAYER	M2 ;
			RECT	0 330.86 0.25 330.96 ;
			LAYER	M3 ;
			RECT	0 330.86 0.25 330.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[99]

	PIN TWENB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 29.18 0.25 29.28 ;
			LAYER	M2 ;
			RECT	0 29.18 0.25 29.28 ;
			LAYER	M3 ;
			RECT	0 29.18 0.25 29.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[9]

	PIN VDDCE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 411.415 21.165 411.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 118.495 21.165 118.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 115.615 21.165 115.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 112.735 21.165 112.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 109.855 21.165 110.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 106.975 21.165 107.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 104.095 21.165 104.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 101.215 21.165 101.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 98.335 21.165 98.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 95.455 21.165 95.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 92.575 21.165 92.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 89.695 21.165 89.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 86.815 21.165 86.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 83.935 21.165 84.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 81.055 21.165 81.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 78.175 21.165 78.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 75.295 21.165 75.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 72.415 21.165 72.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.535 21.165 69.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 66.655 21.165 66.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 63.775 21.165 63.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 60.895 21.165 61.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.015 21.165 58.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.135 21.165 55.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.255 21.165 52.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.375 21.165 49.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 46.495 21.165 46.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 43.615 21.165 43.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 40.735 21.165 40.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 37.855 21.165 38.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 34.975 21.165 35.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.095 21.165 32.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.215 21.165 29.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.335 21.165 26.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.455 21.165 23.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 20.575 21.165 20.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 17.695 21.165 17.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 14.815 21.165 14.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 11.935 21.165 12.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.055 21.165 9.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.175 21.165 6.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.295 21.165 3.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 408.535 21.165 408.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 405.655 21.165 405.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 402.775 21.165 402.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 399.895 21.165 400.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 397.015 21.165 397.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 394.135 21.165 394.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 391.255 21.165 391.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 388.375 21.165 388.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 385.495 21.165 385.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 382.615 21.165 382.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 379.735 21.165 379.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 376.855 21.165 377.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 373.975 21.165 374.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 371.095 21.165 371.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 368.215 21.165 368.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 365.335 21.165 365.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 362.455 21.165 362.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 359.575 21.165 359.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 356.695 21.165 356.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 353.815 21.165 353.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 350.935 21.165 351.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 348.055 21.165 348.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 345.175 21.165 345.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 342.295 21.165 342.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 339.415 21.165 339.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 336.535 21.165 336.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 333.655 21.165 333.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 330.775 21.165 330.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 327.895 21.165 328.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 325.015 21.165 325.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 322.135 21.165 322.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 319.255 21.165 319.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 316.375 21.165 316.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 313.495 21.165 313.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 310.615 21.165 310.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 307.735 21.165 307.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 304.855 21.165 305.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 301.975 21.165 302.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 299.095 21.165 299.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 296.215 21.165 296.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 293.335 21.165 293.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 290.455 21.165 290.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 287.575 21.165 287.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 284.695 21.165 284.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 281.815 21.165 281.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 278.935 21.165 279.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 276.055 21.165 276.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 273.175 21.165 273.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 270.295 21.165 270.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 267.415 21.165 267.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 264.535 21.165 264.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 261.655 21.165 261.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 258.775 21.165 258.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 255.895 21.165 256.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 253.015 21.165 253.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 250.135 21.165 250.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 247.255 21.165 247.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 244.375 21.165 244.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 241.495 21.165 241.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 238.615 21.165 238.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 235.735 21.165 235.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 232.855 21.165 233.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 229.975 21.165 230.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 184.735 21.165 184.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 181.855 21.165 182.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 178.975 21.165 179.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 176.095 21.165 176.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 173.215 21.165 173.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 170.335 21.165 170.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 167.455 21.165 167.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 164.575 21.165 164.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 161.695 21.165 161.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 158.815 21.165 158.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 155.935 21.165 156.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 153.055 21.165 153.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 150.175 21.165 150.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 147.295 21.165 147.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 144.415 21.165 144.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 141.535 21.165 141.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 138.655 21.165 138.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 135.775 21.165 135.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 132.895 21.165 133.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 130.015 21.165 130.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 127.135 21.165 127.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 124.255 21.165 124.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 121.375 21.165 121.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 191.38 21.165 191.57 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 192.36 21.165 192.55 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 195.315 21.165 195.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 199.25 21.165 199.44 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 200.235 21.165 200.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 203.185 21.165 203.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 207.12 21.165 207.31 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 207.615 21.165 207.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 211.55 21.165 211.74 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 214.505 21.165 214.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 215.485 21.165 215.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 219.425 21.165 219.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 222.375 21.165 222.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 223.325 21.165 223.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 414.295 21.165 414.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.415 21.165 0.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 187.095 21.165 187.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 227.615 21.165 227.765 ;
		END

	END VDDCE

	PIN VDDPE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 413.835 21.165 413.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 118.955 21.165 119.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 116.075 21.165 116.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 113.195 21.165 113.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 110.315 21.165 110.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 107.435 21.165 107.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 104.555 21.165 104.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 101.675 21.165 101.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 98.795 21.165 98.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 95.915 21.165 96.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 93.035 21.165 93.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 90.155 21.165 90.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 87.275 21.165 87.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 84.395 21.165 84.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 81.515 21.165 81.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 78.635 21.165 78.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 75.755 21.165 75.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 72.875 21.165 73.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.995 21.165 70.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 67.115 21.165 67.265 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.235 21.165 64.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.355 21.165 61.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.475 21.165 58.625 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.595 21.165 55.745 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.715 21.165 52.865 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.835 21.165 49.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 46.955 21.165 47.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 44.075 21.165 44.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 41.195 21.165 41.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.315 21.165 38.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 35.435 21.165 35.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.555 21.165 32.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.675 21.165 29.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.795 21.165 26.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.915 21.165 24.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 21.035 21.165 21.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 18.155 21.165 18.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.275 21.165 15.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.395 21.165 12.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.515 21.165 9.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.635 21.165 6.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.755 21.165 3.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.875 21.165 1.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 410.955 21.165 411.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 408.075 21.165 408.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 405.195 21.165 405.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 402.315 21.165 402.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 399.435 21.165 399.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 396.555 21.165 396.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 393.675 21.165 393.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 390.795 21.165 390.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 387.915 21.165 388.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 385.035 21.165 385.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 382.155 21.165 382.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 379.275 21.165 379.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 376.395 21.165 376.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 373.515 21.165 373.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 370.635 21.165 370.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 367.755 21.165 367.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 364.875 21.165 365.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 361.995 21.165 362.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 359.115 21.165 359.265 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 356.235 21.165 356.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 353.355 21.165 353.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 350.475 21.165 350.625 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 347.595 21.165 347.745 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 344.715 21.165 344.865 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 341.835 21.165 341.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 338.955 21.165 339.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 336.075 21.165 336.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 333.195 21.165 333.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 330.315 21.165 330.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 327.435 21.165 327.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 324.555 21.165 324.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 321.675 21.165 321.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 318.795 21.165 318.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 315.915 21.165 316.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 313.035 21.165 313.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 310.155 21.165 310.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 307.275 21.165 307.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 304.395 21.165 304.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 301.515 21.165 301.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 298.635 21.165 298.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 295.755 21.165 295.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 292.875 21.165 293.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 289.995 21.165 290.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 287.115 21.165 287.265 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 284.235 21.165 284.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 281.355 21.165 281.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 278.475 21.165 278.625 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 275.595 21.165 275.745 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 272.715 21.165 272.865 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 269.835 21.165 269.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 266.955 21.165 267.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 264.075 21.165 264.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 261.195 21.165 261.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 258.315 21.165 258.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 255.435 21.165 255.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 252.555 21.165 252.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 249.675 21.165 249.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 246.795 21.165 246.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 243.915 21.165 244.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 241.035 21.165 241.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 238.155 21.165 238.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 235.275 21.165 235.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 232.395 21.165 232.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 182.315 21.165 182.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 179.435 21.165 179.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 176.555 21.165 176.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 173.675 21.165 173.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 170.795 21.165 170.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 167.915 21.165 168.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 165.035 21.165 165.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 162.155 21.165 162.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 159.275 21.165 159.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 156.395 21.165 156.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 153.515 21.165 153.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 150.635 21.165 150.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 147.755 21.165 147.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 144.875 21.165 145.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 141.995 21.165 142.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 139.115 21.165 139.265 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 136.235 21.165 136.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 133.355 21.165 133.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 130.475 21.165 130.625 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 127.595 21.165 127.745 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 124.715 21.165 124.865 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 121.835 21.165 121.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 188.425 21.165 188.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 190.43 21.165 190.62 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 193.345 21.165 193.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 194.33 21.165 194.52 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 196.3 21.165 196.49 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 197.28 21.165 197.47 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 198.265 21.165 198.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 201.22 21.165 201.41 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 205.155 21.165 205.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 206.14 21.165 206.33 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 208.6 21.165 208.79 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 209.58 21.165 209.77 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 213.52 21.165 213.71 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 216.47 21.165 216.66 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 217.455 21.165 217.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 218.44 21.165 218.63 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 220.405 21.165 220.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 221.39 21.165 221.58 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 224.31 21.165 224.5 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 226.31 21.165 226.5 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 414.525 21.165 414.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.185 21.165 0.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 186.635 21.165 186.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 228.075 21.165 228.225 ;
		END

	END VDDPE

	PIN VSSE
		USE GROUND ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 414.065 21.165 414.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.645 21.165 0.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 186.865 21.165 187.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 227.845 21.165 227.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 411.185 21.165 411.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 408.305 21.165 408.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 324.785 21.165 324.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 321.905 21.165 322.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 319.025 21.165 319.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 316.145 21.165 316.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 405.425 21.165 405.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 313.265 21.165 313.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 310.385 21.165 310.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 307.505 21.165 307.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 304.625 21.165 304.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 301.745 21.165 301.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 298.865 21.165 299.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 295.985 21.165 296.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 293.105 21.165 293.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 290.225 21.165 290.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 287.345 21.165 287.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 402.545 21.165 402.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 284.465 21.165 284.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 281.585 21.165 281.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 278.705 21.165 278.855 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 275.825 21.165 275.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 272.945 21.165 273.095 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 270.065 21.165 270.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 399.665 21.165 399.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 238.385 21.165 238.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 235.505 21.165 235.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 232.625 21.165 232.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 229.745 21.165 229.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 396.785 21.165 396.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 393.905 21.165 394.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 184.965 21.165 185.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 182.085 21.165 182.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 179.205 21.165 179.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 176.325 21.165 176.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 391.025 21.165 391.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 173.445 21.165 173.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 170.565 21.165 170.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 167.685 21.165 167.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 164.805 21.165 164.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 161.925 21.165 162.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 159.045 21.165 159.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 156.165 21.165 156.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 153.285 21.165 153.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 150.405 21.165 150.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 147.525 21.165 147.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 388.145 21.165 388.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 144.645 21.165 144.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 141.765 21.165 141.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 138.885 21.165 139.035 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 136.005 21.165 136.155 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 133.125 21.165 133.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 130.245 21.165 130.395 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 127.365 21.165 127.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 124.485 21.165 124.635 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 121.605 21.165 121.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 118.725 21.165 118.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 385.265 21.165 385.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 115.845 21.165 115.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 112.965 21.165 113.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 110.085 21.165 110.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 107.205 21.165 107.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 104.325 21.165 104.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 101.445 21.165 101.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 98.565 21.165 98.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 95.685 21.165 95.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 92.805 21.165 92.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 89.925 21.165 90.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 382.385 21.165 382.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 87.045 21.165 87.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 84.165 21.165 84.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 81.285 21.165 81.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 78.405 21.165 78.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 75.525 21.165 75.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 72.645 21.165 72.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.765 21.165 69.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 66.885 21.165 67.035 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 379.505 21.165 379.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 376.625 21.165 376.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.685 21.165 23.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 20.805 21.165 20.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 17.925 21.165 18.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.045 21.165 15.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.165 21.165 12.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.285 21.165 9.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.405 21.165 6.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.525 21.165 3.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 373.745 21.165 373.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 370.865 21.165 371.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 367.985 21.165 368.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 413.605 21.165 413.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 344.485 21.165 344.635 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 341.605 21.165 341.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 338.725 21.165 338.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 335.845 21.165 335.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 332.965 21.165 333.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 407.845 21.165 407.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 330.085 21.165 330.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 327.205 21.165 327.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 324.325 21.165 324.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 321.445 21.165 321.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 318.565 21.165 318.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 315.685 21.165 315.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 312.805 21.165 312.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 309.925 21.165 310.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 307.045 21.165 307.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 304.165 21.165 304.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 404.965 21.165 405.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 301.285 21.165 301.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 298.405 21.165 298.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 295.525 21.165 295.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 292.645 21.165 292.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 289.765 21.165 289.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 286.885 21.165 287.035 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 284.005 21.165 284.155 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 281.125 21.165 281.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 278.245 21.165 278.395 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 275.365 21.165 275.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 402.085 21.165 402.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 272.485 21.165 272.635 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 269.605 21.165 269.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 266.725 21.165 266.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 263.845 21.165 263.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 260.965 21.165 261.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 258.085 21.165 258.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 255.205 21.165 255.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 252.325 21.165 252.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 249.445 21.165 249.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 246.565 21.165 246.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 399.205 21.165 399.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 243.685 21.165 243.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 240.805 21.165 240.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 237.925 21.165 238.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 235.045 21.165 235.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 232.165 21.165 232.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 396.325 21.165 396.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 393.445 21.165 393.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 182.545 21.165 182.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 179.665 21.165 179.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 176.785 21.165 176.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 173.905 21.165 174.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 171.025 21.165 171.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 168.145 21.165 168.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 165.265 21.165 165.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 162.385 21.165 162.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 159.505 21.165 159.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 390.565 21.165 390.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 156.625 21.165 156.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 153.745 21.165 153.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 150.865 21.165 151.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 147.985 21.165 148.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 145.105 21.165 145.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 142.225 21.165 142.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 139.345 21.165 139.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 136.465 21.165 136.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 133.585 21.165 133.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 130.705 21.165 130.855 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 387.685 21.165 387.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 127.825 21.165 127.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 124.945 21.165 125.095 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 122.065 21.165 122.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 119.185 21.165 119.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 116.305 21.165 116.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 113.425 21.165 113.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 110.545 21.165 110.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 107.665 21.165 107.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 104.785 21.165 104.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 101.905 21.165 102.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 384.805 21.165 384.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 99.025 21.165 99.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 96.145 21.165 96.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 93.265 21.165 93.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 90.385 21.165 90.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 87.505 21.165 87.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 84.625 21.165 84.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 81.745 21.165 81.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 78.865 21.165 79.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 75.985 21.165 76.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 73.105 21.165 73.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 381.925 21.165 382.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 70.225 21.165 70.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 67.345 21.165 67.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.825 21.165 55.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.945 21.165 53.095 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 50.065 21.165 50.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 47.185 21.165 47.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 44.305 21.165 44.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 379.045 21.165 379.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 41.425 21.165 41.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.545 21.165 38.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 35.665 21.165 35.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.785 21.165 32.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.905 21.165 30.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 27.025 21.165 27.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 24.145 21.165 24.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 21.265 21.165 21.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 18.385 21.165 18.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.505 21.165 15.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 376.165 21.165 376.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.625 21.165 12.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.745 21.165 9.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.865 21.165 7.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.985 21.165 4.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 1.105 21.165 1.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 373.285 21.165 373.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 370.405 21.165 370.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 367.525 21.165 367.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 410.725 21.165 410.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 356.005 21.165 356.155 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 353.125 21.165 353.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 350.245 21.165 350.395 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 347.365 21.165 347.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 187.935 21.165 188.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 188.915 21.165 189.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 190.885 21.165 191.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 191.87 21.165 192.06 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 194.825 21.165 195.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 195.805 21.165 195.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 196.79 21.165 196.98 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 198.76 21.165 198.95 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 199.73 21.165 199.94 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 200.725 21.165 200.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 202.7 21.165 202.89 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 203.68 21.165 203.87 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 206.63 21.165 206.82 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 208.105 21.165 208.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 211.055 21.165 211.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 212.045 21.165 212.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 214.01 21.165 214.2 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 214.985 21.165 215.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 215.98 21.165 216.17 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 217.945 21.165 218.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 218.93 21.165 219.12 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 219.915 21.165 220.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 222.855 21.165 223.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 223.85 21.165 224.04 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 225.82 21.165 226.01 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 226.805 21.165 226.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.005 21.165 64.155 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.125 21.165 61.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.245 21.165 58.395 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.365 21.165 55.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.485 21.165 52.635 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.605 21.165 49.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 46.725 21.165 46.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 43.845 21.165 43.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 40.965 21.165 41.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.085 21.165 38.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 35.205 21.165 35.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.325 21.165 32.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.445 21.165 29.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.565 21.165 26.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 365.105 21.165 365.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 362.225 21.165 362.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 359.345 21.165 359.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 356.465 21.165 356.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 353.585 21.165 353.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 350.705 21.165 350.855 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 347.825 21.165 347.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 344.945 21.165 345.095 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 342.065 21.165 342.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 339.185 21.165 339.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 336.305 21.165 336.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 333.425 21.165 333.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 330.545 21.165 330.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 327.665 21.165 327.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 267.185 21.165 267.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 264.305 21.165 264.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 261.425 21.165 261.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 258.545 21.165 258.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 255.665 21.165 255.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 252.785 21.165 252.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 249.905 21.165 250.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 247.025 21.165 247.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 244.145 21.165 244.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 241.265 21.165 241.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.465 21.165 64.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.585 21.165 61.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.705 21.165 58.855 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 364.645 21.165 364.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 361.765 21.165 361.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 358.885 21.165 359.035 ;
		END

	END VSSE

	PIN WENB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 1.995 0.25 2.095 ;
			LAYER	M2 ;
			RECT	0 1.995 0.25 2.095 ;
			LAYER	M3 ;
			RECT	0 1.995 0.25 2.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[0]

	PIN WENB[100]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 335.005 0.25 335.105 ;
			LAYER	M2 ;
			RECT	0 335.005 0.25 335.105 ;
			LAYER	M3 ;
			RECT	0 335.005 0.25 335.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[100]

	PIN WENB[101]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 337.885 0.25 337.985 ;
			LAYER	M2 ;
			RECT	0 337.885 0.25 337.985 ;
			LAYER	M3 ;
			RECT	0 337.885 0.25 337.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[101]

	PIN WENB[102]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 340.765 0.25 340.865 ;
			LAYER	M2 ;
			RECT	0 340.765 0.25 340.865 ;
			LAYER	M3 ;
			RECT	0 340.765 0.25 340.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[102]

	PIN WENB[103]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 343.645 0.25 343.745 ;
			LAYER	M2 ;
			RECT	0 343.645 0.25 343.745 ;
			LAYER	M3 ;
			RECT	0 343.645 0.25 343.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[103]

	PIN WENB[104]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 346.525 0.25 346.625 ;
			LAYER	M2 ;
			RECT	0 346.525 0.25 346.625 ;
			LAYER	M3 ;
			RECT	0 346.525 0.25 346.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[104]

	PIN WENB[105]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 349.405 0.25 349.505 ;
			LAYER	M2 ;
			RECT	0 349.405 0.25 349.505 ;
			LAYER	M3 ;
			RECT	0 349.405 0.25 349.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[105]

	PIN WENB[106]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 352.285 0.25 352.385 ;
			LAYER	M2 ;
			RECT	0 352.285 0.25 352.385 ;
			LAYER	M3 ;
			RECT	0 352.285 0.25 352.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[106]

	PIN WENB[107]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 355.165 0.25 355.265 ;
			LAYER	M2 ;
			RECT	0 355.165 0.25 355.265 ;
			LAYER	M3 ;
			RECT	0 355.165 0.25 355.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[107]

	PIN WENB[108]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 358.045 0.25 358.145 ;
			LAYER	M2 ;
			RECT	0 358.045 0.25 358.145 ;
			LAYER	M3 ;
			RECT	0 358.045 0.25 358.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[108]

	PIN WENB[109]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 360.925 0.25 361.025 ;
			LAYER	M2 ;
			RECT	0 360.925 0.25 361.025 ;
			LAYER	M3 ;
			RECT	0 360.925 0.25 361.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[109]

	PIN WENB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.795 0.25 30.895 ;
			LAYER	M2 ;
			RECT	0 30.795 0.25 30.895 ;
			LAYER	M3 ;
			RECT	0 30.795 0.25 30.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[10]

	PIN WENB[110]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 363.805 0.25 363.905 ;
			LAYER	M2 ;
			RECT	0 363.805 0.25 363.905 ;
			LAYER	M3 ;
			RECT	0 363.805 0.25 363.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[110]

	PIN WENB[111]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 366.685 0.25 366.785 ;
			LAYER	M2 ;
			RECT	0 366.685 0.25 366.785 ;
			LAYER	M3 ;
			RECT	0 366.685 0.25 366.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[111]

	PIN WENB[112]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 369.565 0.25 369.665 ;
			LAYER	M2 ;
			RECT	0 369.565 0.25 369.665 ;
			LAYER	M3 ;
			RECT	0 369.565 0.25 369.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[112]

	PIN WENB[113]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 372.445 0.25 372.545 ;
			LAYER	M2 ;
			RECT	0 372.445 0.25 372.545 ;
			LAYER	M3 ;
			RECT	0 372.445 0.25 372.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[113]

	PIN WENB[114]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 375.325 0.25 375.425 ;
			LAYER	M2 ;
			RECT	0 375.325 0.25 375.425 ;
			LAYER	M3 ;
			RECT	0 375.325 0.25 375.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[114]

	PIN WENB[115]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 378.205 0.25 378.305 ;
			LAYER	M2 ;
			RECT	0 378.205 0.25 378.305 ;
			LAYER	M3 ;
			RECT	0 378.205 0.25 378.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[115]

	PIN WENB[116]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 381.085 0.25 381.185 ;
			LAYER	M2 ;
			RECT	0 381.085 0.25 381.185 ;
			LAYER	M3 ;
			RECT	0 381.085 0.25 381.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[116]

	PIN WENB[117]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 383.965 0.25 384.065 ;
			LAYER	M2 ;
			RECT	0 383.965 0.25 384.065 ;
			LAYER	M3 ;
			RECT	0 383.965 0.25 384.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[117]

	PIN WENB[118]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 386.845 0.25 386.945 ;
			LAYER	M2 ;
			RECT	0 386.845 0.25 386.945 ;
			LAYER	M3 ;
			RECT	0 386.845 0.25 386.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[118]

	PIN WENB[119]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 389.725 0.25 389.825 ;
			LAYER	M2 ;
			RECT	0 389.725 0.25 389.825 ;
			LAYER	M3 ;
			RECT	0 389.725 0.25 389.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[119]

	PIN WENB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.675 0.25 33.775 ;
			LAYER	M2 ;
			RECT	0 33.675 0.25 33.775 ;
			LAYER	M3 ;
			RECT	0 33.675 0.25 33.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[11]

	PIN WENB[120]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 392.605 0.25 392.705 ;
			LAYER	M2 ;
			RECT	0 392.605 0.25 392.705 ;
			LAYER	M3 ;
			RECT	0 392.605 0.25 392.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[120]

	PIN WENB[121]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 395.485 0.25 395.585 ;
			LAYER	M2 ;
			RECT	0 395.485 0.25 395.585 ;
			LAYER	M3 ;
			RECT	0 395.485 0.25 395.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[121]

	PIN WENB[122]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 398.365 0.25 398.465 ;
			LAYER	M2 ;
			RECT	0 398.365 0.25 398.465 ;
			LAYER	M3 ;
			RECT	0 398.365 0.25 398.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[122]

	PIN WENB[123]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 401.245 0.25 401.345 ;
			LAYER	M2 ;
			RECT	0 401.245 0.25 401.345 ;
			LAYER	M3 ;
			RECT	0 401.245 0.25 401.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[123]

	PIN WENB[124]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 404.125 0.25 404.225 ;
			LAYER	M2 ;
			RECT	0 404.125 0.25 404.225 ;
			LAYER	M3 ;
			RECT	0 404.125 0.25 404.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[124]

	PIN WENB[125]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 407.005 0.25 407.105 ;
			LAYER	M2 ;
			RECT	0 407.005 0.25 407.105 ;
			LAYER	M3 ;
			RECT	0 407.005 0.25 407.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[125]

	PIN WENB[126]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 409.885 0.25 409.985 ;
			LAYER	M2 ;
			RECT	0 409.885 0.25 409.985 ;
			LAYER	M3 ;
			RECT	0 409.885 0.25 409.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[126]

	PIN WENB[127]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 412.765 0.25 412.865 ;
			LAYER	M2 ;
			RECT	0 412.765 0.25 412.865 ;
			LAYER	M3 ;
			RECT	0 412.765 0.25 412.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[127]

	PIN WENB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.555 0.25 36.655 ;
			LAYER	M2 ;
			RECT	0 36.555 0.25 36.655 ;
			LAYER	M3 ;
			RECT	0 36.555 0.25 36.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[12]

	PIN WENB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.435 0.25 39.535 ;
			LAYER	M2 ;
			RECT	0 39.435 0.25 39.535 ;
			LAYER	M3 ;
			RECT	0 39.435 0.25 39.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[13]

	PIN WENB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.315 0.25 42.415 ;
			LAYER	M2 ;
			RECT	0 42.315 0.25 42.415 ;
			LAYER	M3 ;
			RECT	0 42.315 0.25 42.415 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[14]

	PIN WENB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 45.195 0.25 45.295 ;
			LAYER	M2 ;
			RECT	0 45.195 0.25 45.295 ;
			LAYER	M3 ;
			RECT	0 45.195 0.25 45.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[15]

	PIN WENB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 48.075 0.25 48.175 ;
			LAYER	M2 ;
			RECT	0 48.075 0.25 48.175 ;
			LAYER	M3 ;
			RECT	0 48.075 0.25 48.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[16]

	PIN WENB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 50.955 0.25 51.055 ;
			LAYER	M2 ;
			RECT	0 50.955 0.25 51.055 ;
			LAYER	M3 ;
			RECT	0 50.955 0.25 51.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[17]

	PIN WENB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 53.835 0.25 53.935 ;
			LAYER	M2 ;
			RECT	0 53.835 0.25 53.935 ;
			LAYER	M3 ;
			RECT	0 53.835 0.25 53.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[18]

	PIN WENB[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.715 0.25 56.815 ;
			LAYER	M2 ;
			RECT	0 56.715 0.25 56.815 ;
			LAYER	M3 ;
			RECT	0 56.715 0.25 56.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[19]

	PIN WENB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 4.875 0.25 4.975 ;
			LAYER	M2 ;
			RECT	0 4.875 0.25 4.975 ;
			LAYER	M3 ;
			RECT	0 4.875 0.25 4.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[1]

	PIN WENB[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.595 0.25 59.695 ;
			LAYER	M2 ;
			RECT	0 59.595 0.25 59.695 ;
			LAYER	M3 ;
			RECT	0 59.595 0.25 59.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[20]

	PIN WENB[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.475 0.25 62.575 ;
			LAYER	M2 ;
			RECT	0 62.475 0.25 62.575 ;
			LAYER	M3 ;
			RECT	0 62.475 0.25 62.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[21]

	PIN WENB[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.355 0.25 65.455 ;
			LAYER	M2 ;
			RECT	0 65.355 0.25 65.455 ;
			LAYER	M3 ;
			RECT	0 65.355 0.25 65.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[22]

	PIN WENB[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 68.235 0.25 68.335 ;
			LAYER	M2 ;
			RECT	0 68.235 0.25 68.335 ;
			LAYER	M3 ;
			RECT	0 68.235 0.25 68.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[23]

	PIN WENB[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 71.115 0.25 71.215 ;
			LAYER	M2 ;
			RECT	0 71.115 0.25 71.215 ;
			LAYER	M3 ;
			RECT	0 71.115 0.25 71.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[24]

	PIN WENB[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 73.995 0.25 74.095 ;
			LAYER	M2 ;
			RECT	0 73.995 0.25 74.095 ;
			LAYER	M3 ;
			RECT	0 73.995 0.25 74.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[25]

	PIN WENB[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 76.875 0.25 76.975 ;
			LAYER	M2 ;
			RECT	0 76.875 0.25 76.975 ;
			LAYER	M3 ;
			RECT	0 76.875 0.25 76.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[26]

	PIN WENB[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.755 0.25 79.855 ;
			LAYER	M2 ;
			RECT	0 79.755 0.25 79.855 ;
			LAYER	M3 ;
			RECT	0 79.755 0.25 79.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[27]

	PIN WENB[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.635 0.25 82.735 ;
			LAYER	M2 ;
			RECT	0 82.635 0.25 82.735 ;
			LAYER	M3 ;
			RECT	0 82.635 0.25 82.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[28]

	PIN WENB[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 85.515 0.25 85.615 ;
			LAYER	M2 ;
			RECT	0 85.515 0.25 85.615 ;
			LAYER	M3 ;
			RECT	0 85.515 0.25 85.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[29]

	PIN WENB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.755 0.25 7.855 ;
			LAYER	M2 ;
			RECT	0 7.755 0.25 7.855 ;
			LAYER	M3 ;
			RECT	0 7.755 0.25 7.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[2]

	PIN WENB[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 88.395 0.25 88.495 ;
			LAYER	M2 ;
			RECT	0 88.395 0.25 88.495 ;
			LAYER	M3 ;
			RECT	0 88.395 0.25 88.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[30]

	PIN WENB[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 91.275 0.25 91.375 ;
			LAYER	M2 ;
			RECT	0 91.275 0.25 91.375 ;
			LAYER	M3 ;
			RECT	0 91.275 0.25 91.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[31]

	PIN WENB[32]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 94.155 0.25 94.255 ;
			LAYER	M2 ;
			RECT	0 94.155 0.25 94.255 ;
			LAYER	M3 ;
			RECT	0 94.155 0.25 94.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[32]

	PIN WENB[33]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 97.035 0.25 97.135 ;
			LAYER	M2 ;
			RECT	0 97.035 0.25 97.135 ;
			LAYER	M3 ;
			RECT	0 97.035 0.25 97.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[33]

	PIN WENB[34]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 99.915 0.25 100.015 ;
			LAYER	M2 ;
			RECT	0 99.915 0.25 100.015 ;
			LAYER	M3 ;
			RECT	0 99.915 0.25 100.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[34]

	PIN WENB[35]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 102.795 0.25 102.895 ;
			LAYER	M2 ;
			RECT	0 102.795 0.25 102.895 ;
			LAYER	M3 ;
			RECT	0 102.795 0.25 102.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[35]

	PIN WENB[36]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 105.675 0.25 105.775 ;
			LAYER	M2 ;
			RECT	0 105.675 0.25 105.775 ;
			LAYER	M3 ;
			RECT	0 105.675 0.25 105.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[36]

	PIN WENB[37]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 108.555 0.25 108.655 ;
			LAYER	M2 ;
			RECT	0 108.555 0.25 108.655 ;
			LAYER	M3 ;
			RECT	0 108.555 0.25 108.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[37]

	PIN WENB[38]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 111.435 0.25 111.535 ;
			LAYER	M2 ;
			RECT	0 111.435 0.25 111.535 ;
			LAYER	M3 ;
			RECT	0 111.435 0.25 111.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[38]

	PIN WENB[39]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 114.315 0.25 114.415 ;
			LAYER	M2 ;
			RECT	0 114.315 0.25 114.415 ;
			LAYER	M3 ;
			RECT	0 114.315 0.25 114.415 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[39]

	PIN WENB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.635 0.25 10.735 ;
			LAYER	M2 ;
			RECT	0 10.635 0.25 10.735 ;
			LAYER	M3 ;
			RECT	0 10.635 0.25 10.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[3]

	PIN WENB[40]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 117.195 0.25 117.295 ;
			LAYER	M2 ;
			RECT	0 117.195 0.25 117.295 ;
			LAYER	M3 ;
			RECT	0 117.195 0.25 117.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[40]

	PIN WENB[41]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 120.075 0.25 120.175 ;
			LAYER	M2 ;
			RECT	0 120.075 0.25 120.175 ;
			LAYER	M3 ;
			RECT	0 120.075 0.25 120.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[41]

	PIN WENB[42]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 122.955 0.25 123.055 ;
			LAYER	M2 ;
			RECT	0 122.955 0.25 123.055 ;
			LAYER	M3 ;
			RECT	0 122.955 0.25 123.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[42]

	PIN WENB[43]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 125.835 0.25 125.935 ;
			LAYER	M2 ;
			RECT	0 125.835 0.25 125.935 ;
			LAYER	M3 ;
			RECT	0 125.835 0.25 125.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[43]

	PIN WENB[44]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 128.715 0.25 128.815 ;
			LAYER	M2 ;
			RECT	0 128.715 0.25 128.815 ;
			LAYER	M3 ;
			RECT	0 128.715 0.25 128.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[44]

	PIN WENB[45]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 131.595 0.25 131.695 ;
			LAYER	M2 ;
			RECT	0 131.595 0.25 131.695 ;
			LAYER	M3 ;
			RECT	0 131.595 0.25 131.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[45]

	PIN WENB[46]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 134.475 0.25 134.575 ;
			LAYER	M2 ;
			RECT	0 134.475 0.25 134.575 ;
			LAYER	M3 ;
			RECT	0 134.475 0.25 134.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[46]

	PIN WENB[47]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 137.355 0.25 137.455 ;
			LAYER	M2 ;
			RECT	0 137.355 0.25 137.455 ;
			LAYER	M3 ;
			RECT	0 137.355 0.25 137.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[47]

	PIN WENB[48]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 140.235 0.25 140.335 ;
			LAYER	M2 ;
			RECT	0 140.235 0.25 140.335 ;
			LAYER	M3 ;
			RECT	0 140.235 0.25 140.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[48]

	PIN WENB[49]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 143.115 0.25 143.215 ;
			LAYER	M2 ;
			RECT	0 143.115 0.25 143.215 ;
			LAYER	M3 ;
			RECT	0 143.115 0.25 143.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[49]

	PIN WENB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.515 0.25 13.615 ;
			LAYER	M2 ;
			RECT	0 13.515 0.25 13.615 ;
			LAYER	M3 ;
			RECT	0 13.515 0.25 13.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[4]

	PIN WENB[50]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 145.995 0.25 146.095 ;
			LAYER	M2 ;
			RECT	0 145.995 0.25 146.095 ;
			LAYER	M3 ;
			RECT	0 145.995 0.25 146.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[50]

	PIN WENB[51]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 148.875 0.25 148.975 ;
			LAYER	M2 ;
			RECT	0 148.875 0.25 148.975 ;
			LAYER	M3 ;
			RECT	0 148.875 0.25 148.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[51]

	PIN WENB[52]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 151.755 0.25 151.855 ;
			LAYER	M2 ;
			RECT	0 151.755 0.25 151.855 ;
			LAYER	M3 ;
			RECT	0 151.755 0.25 151.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[52]

	PIN WENB[53]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 154.635 0.25 154.735 ;
			LAYER	M2 ;
			RECT	0 154.635 0.25 154.735 ;
			LAYER	M3 ;
			RECT	0 154.635 0.25 154.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[53]

	PIN WENB[54]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 157.515 0.25 157.615 ;
			LAYER	M2 ;
			RECT	0 157.515 0.25 157.615 ;
			LAYER	M3 ;
			RECT	0 157.515 0.25 157.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[54]

	PIN WENB[55]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 160.395 0.25 160.495 ;
			LAYER	M2 ;
			RECT	0 160.395 0.25 160.495 ;
			LAYER	M3 ;
			RECT	0 160.395 0.25 160.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[55]

	PIN WENB[56]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 163.275 0.25 163.375 ;
			LAYER	M2 ;
			RECT	0 163.275 0.25 163.375 ;
			LAYER	M3 ;
			RECT	0 163.275 0.25 163.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[56]

	PIN WENB[57]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 166.155 0.25 166.255 ;
			LAYER	M2 ;
			RECT	0 166.155 0.25 166.255 ;
			LAYER	M3 ;
			RECT	0 166.155 0.25 166.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[57]

	PIN WENB[58]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 169.035 0.25 169.135 ;
			LAYER	M2 ;
			RECT	0 169.035 0.25 169.135 ;
			LAYER	M3 ;
			RECT	0 169.035 0.25 169.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[58]

	PIN WENB[59]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 171.915 0.25 172.015 ;
			LAYER	M2 ;
			RECT	0 171.915 0.25 172.015 ;
			LAYER	M3 ;
			RECT	0 171.915 0.25 172.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[59]

	PIN WENB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.395 0.25 16.495 ;
			LAYER	M2 ;
			RECT	0 16.395 0.25 16.495 ;
			LAYER	M3 ;
			RECT	0 16.395 0.25 16.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[5]

	PIN WENB[60]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 174.795 0.25 174.895 ;
			LAYER	M2 ;
			RECT	0 174.795 0.25 174.895 ;
			LAYER	M3 ;
			RECT	0 174.795 0.25 174.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[60]

	PIN WENB[61]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 177.675 0.25 177.775 ;
			LAYER	M2 ;
			RECT	0 177.675 0.25 177.775 ;
			LAYER	M3 ;
			RECT	0 177.675 0.25 177.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[61]

	PIN WENB[62]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 180.555 0.25 180.655 ;
			LAYER	M2 ;
			RECT	0 180.555 0.25 180.655 ;
			LAYER	M3 ;
			RECT	0 180.555 0.25 180.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[62]

	PIN WENB[63]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 183.435 0.25 183.535 ;
			LAYER	M2 ;
			RECT	0 183.435 0.25 183.535 ;
			LAYER	M3 ;
			RECT	0 183.435 0.25 183.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[63]

	PIN WENB[64]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 231.325 0.25 231.425 ;
			LAYER	M2 ;
			RECT	0 231.325 0.25 231.425 ;
			LAYER	M3 ;
			RECT	0 231.325 0.25 231.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[64]

	PIN WENB[65]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 234.205 0.25 234.305 ;
			LAYER	M2 ;
			RECT	0 234.205 0.25 234.305 ;
			LAYER	M3 ;
			RECT	0 234.205 0.25 234.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[65]

	PIN WENB[66]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 237.085 0.25 237.185 ;
			LAYER	M2 ;
			RECT	0 237.085 0.25 237.185 ;
			LAYER	M3 ;
			RECT	0 237.085 0.25 237.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[66]

	PIN WENB[67]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 239.965 0.25 240.065 ;
			LAYER	M2 ;
			RECT	0 239.965 0.25 240.065 ;
			LAYER	M3 ;
			RECT	0 239.965 0.25 240.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[67]

	PIN WENB[68]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 242.845 0.25 242.945 ;
			LAYER	M2 ;
			RECT	0 242.845 0.25 242.945 ;
			LAYER	M3 ;
			RECT	0 242.845 0.25 242.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[68]

	PIN WENB[69]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 245.725 0.25 245.825 ;
			LAYER	M2 ;
			RECT	0 245.725 0.25 245.825 ;
			LAYER	M3 ;
			RECT	0 245.725 0.25 245.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[69]

	PIN WENB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.275 0.25 19.375 ;
			LAYER	M2 ;
			RECT	0 19.275 0.25 19.375 ;
			LAYER	M3 ;
			RECT	0 19.275 0.25 19.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[6]

	PIN WENB[70]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 248.605 0.25 248.705 ;
			LAYER	M2 ;
			RECT	0 248.605 0.25 248.705 ;
			LAYER	M3 ;
			RECT	0 248.605 0.25 248.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[70]

	PIN WENB[71]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 251.485 0.25 251.585 ;
			LAYER	M2 ;
			RECT	0 251.485 0.25 251.585 ;
			LAYER	M3 ;
			RECT	0 251.485 0.25 251.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[71]

	PIN WENB[72]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 254.365 0.25 254.465 ;
			LAYER	M2 ;
			RECT	0 254.365 0.25 254.465 ;
			LAYER	M3 ;
			RECT	0 254.365 0.25 254.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[72]

	PIN WENB[73]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 257.245 0.25 257.345 ;
			LAYER	M2 ;
			RECT	0 257.245 0.25 257.345 ;
			LAYER	M3 ;
			RECT	0 257.245 0.25 257.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[73]

	PIN WENB[74]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 260.125 0.25 260.225 ;
			LAYER	M2 ;
			RECT	0 260.125 0.25 260.225 ;
			LAYER	M3 ;
			RECT	0 260.125 0.25 260.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[74]

	PIN WENB[75]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 263.005 0.25 263.105 ;
			LAYER	M2 ;
			RECT	0 263.005 0.25 263.105 ;
			LAYER	M3 ;
			RECT	0 263.005 0.25 263.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[75]

	PIN WENB[76]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 265.885 0.25 265.985 ;
			LAYER	M2 ;
			RECT	0 265.885 0.25 265.985 ;
			LAYER	M3 ;
			RECT	0 265.885 0.25 265.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[76]

	PIN WENB[77]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 268.765 0.25 268.865 ;
			LAYER	M2 ;
			RECT	0 268.765 0.25 268.865 ;
			LAYER	M3 ;
			RECT	0 268.765 0.25 268.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[77]

	PIN WENB[78]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 271.645 0.25 271.745 ;
			LAYER	M2 ;
			RECT	0 271.645 0.25 271.745 ;
			LAYER	M3 ;
			RECT	0 271.645 0.25 271.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[78]

	PIN WENB[79]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 274.525 0.25 274.625 ;
			LAYER	M2 ;
			RECT	0 274.525 0.25 274.625 ;
			LAYER	M3 ;
			RECT	0 274.525 0.25 274.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[79]

	PIN WENB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.155 0.25 22.255 ;
			LAYER	M2 ;
			RECT	0 22.155 0.25 22.255 ;
			LAYER	M3 ;
			RECT	0 22.155 0.25 22.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[7]

	PIN WENB[80]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 277.405 0.25 277.505 ;
			LAYER	M2 ;
			RECT	0 277.405 0.25 277.505 ;
			LAYER	M3 ;
			RECT	0 277.405 0.25 277.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[80]

	PIN WENB[81]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 280.285 0.25 280.385 ;
			LAYER	M2 ;
			RECT	0 280.285 0.25 280.385 ;
			LAYER	M3 ;
			RECT	0 280.285 0.25 280.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[81]

	PIN WENB[82]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 283.165 0.25 283.265 ;
			LAYER	M2 ;
			RECT	0 283.165 0.25 283.265 ;
			LAYER	M3 ;
			RECT	0 283.165 0.25 283.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[82]

	PIN WENB[83]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 286.045 0.25 286.145 ;
			LAYER	M2 ;
			RECT	0 286.045 0.25 286.145 ;
			LAYER	M3 ;
			RECT	0 286.045 0.25 286.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[83]

	PIN WENB[84]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 288.925 0.25 289.025 ;
			LAYER	M2 ;
			RECT	0 288.925 0.25 289.025 ;
			LAYER	M3 ;
			RECT	0 288.925 0.25 289.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[84]

	PIN WENB[85]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 291.805 0.25 291.905 ;
			LAYER	M2 ;
			RECT	0 291.805 0.25 291.905 ;
			LAYER	M3 ;
			RECT	0 291.805 0.25 291.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[85]

	PIN WENB[86]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 294.685 0.25 294.785 ;
			LAYER	M2 ;
			RECT	0 294.685 0.25 294.785 ;
			LAYER	M3 ;
			RECT	0 294.685 0.25 294.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[86]

	PIN WENB[87]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 297.565 0.25 297.665 ;
			LAYER	M2 ;
			RECT	0 297.565 0.25 297.665 ;
			LAYER	M3 ;
			RECT	0 297.565 0.25 297.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[87]

	PIN WENB[88]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 300.445 0.25 300.545 ;
			LAYER	M2 ;
			RECT	0 300.445 0.25 300.545 ;
			LAYER	M3 ;
			RECT	0 300.445 0.25 300.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[88]

	PIN WENB[89]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 303.325 0.25 303.425 ;
			LAYER	M2 ;
			RECT	0 303.325 0.25 303.425 ;
			LAYER	M3 ;
			RECT	0 303.325 0.25 303.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[89]

	PIN WENB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.035 0.25 25.135 ;
			LAYER	M2 ;
			RECT	0 25.035 0.25 25.135 ;
			LAYER	M3 ;
			RECT	0 25.035 0.25 25.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[8]

	PIN WENB[90]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 306.205 0.25 306.305 ;
			LAYER	M2 ;
			RECT	0 306.205 0.25 306.305 ;
			LAYER	M3 ;
			RECT	0 306.205 0.25 306.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[90]

	PIN WENB[91]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 309.085 0.25 309.185 ;
			LAYER	M2 ;
			RECT	0 309.085 0.25 309.185 ;
			LAYER	M3 ;
			RECT	0 309.085 0.25 309.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[91]

	PIN WENB[92]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 311.965 0.25 312.065 ;
			LAYER	M2 ;
			RECT	0 311.965 0.25 312.065 ;
			LAYER	M3 ;
			RECT	0 311.965 0.25 312.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[92]

	PIN WENB[93]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 314.845 0.25 314.945 ;
			LAYER	M2 ;
			RECT	0 314.845 0.25 314.945 ;
			LAYER	M3 ;
			RECT	0 314.845 0.25 314.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[93]

	PIN WENB[94]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 317.725 0.25 317.825 ;
			LAYER	M2 ;
			RECT	0 317.725 0.25 317.825 ;
			LAYER	M3 ;
			RECT	0 317.725 0.25 317.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[94]

	PIN WENB[95]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 320.605 0.25 320.705 ;
			LAYER	M2 ;
			RECT	0 320.605 0.25 320.705 ;
			LAYER	M3 ;
			RECT	0 320.605 0.25 320.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[95]

	PIN WENB[96]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 323.485 0.25 323.585 ;
			LAYER	M2 ;
			RECT	0 323.485 0.25 323.585 ;
			LAYER	M3 ;
			RECT	0 323.485 0.25 323.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[96]

	PIN WENB[97]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 326.365 0.25 326.465 ;
			LAYER	M2 ;
			RECT	0 326.365 0.25 326.465 ;
			LAYER	M3 ;
			RECT	0 326.365 0.25 326.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[97]

	PIN WENB[98]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 329.245 0.25 329.345 ;
			LAYER	M2 ;
			RECT	0 329.245 0.25 329.345 ;
			LAYER	M3 ;
			RECT	0 329.245 0.25 329.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[98]

	PIN WENB[99]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 332.125 0.25 332.225 ;
			LAYER	M2 ;
			RECT	0 332.125 0.25 332.225 ;
			LAYER	M3 ;
			RECT	0 332.125 0.25 332.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[99]

	PIN WENB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 27.915 0.25 28.015 ;
			LAYER	M2 ;
			RECT	0 27.915 0.25 28.015 ;
			LAYER	M3 ;
			RECT	0 27.915 0.25 28.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[9]

	PIN WENYB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 1.73 0.25 1.83 ;
			LAYER	M2 ;
			RECT	0 1.73 0.25 1.83 ;
			LAYER	M3 ;
			RECT	0 1.73 0.25 1.83 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[0]

	PIN WENYB[100]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 335.27 0.25 335.37 ;
			LAYER	M2 ;
			RECT	0 335.27 0.25 335.37 ;
			LAYER	M3 ;
			RECT	0 335.27 0.25 335.37 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[100]

	PIN WENYB[101]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 338.15 0.25 338.25 ;
			LAYER	M2 ;
			RECT	0 338.15 0.25 338.25 ;
			LAYER	M3 ;
			RECT	0 338.15 0.25 338.25 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[101]

	PIN WENYB[102]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 341.03 0.25 341.13 ;
			LAYER	M2 ;
			RECT	0 341.03 0.25 341.13 ;
			LAYER	M3 ;
			RECT	0 341.03 0.25 341.13 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[102]

	PIN WENYB[103]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 343.91 0.25 344.01 ;
			LAYER	M2 ;
			RECT	0 343.91 0.25 344.01 ;
			LAYER	M3 ;
			RECT	0 343.91 0.25 344.01 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[103]

	PIN WENYB[104]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 346.79 0.25 346.89 ;
			LAYER	M2 ;
			RECT	0 346.79 0.25 346.89 ;
			LAYER	M3 ;
			RECT	0 346.79 0.25 346.89 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[104]

	PIN WENYB[105]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 349.67 0.25 349.77 ;
			LAYER	M2 ;
			RECT	0 349.67 0.25 349.77 ;
			LAYER	M3 ;
			RECT	0 349.67 0.25 349.77 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[105]

	PIN WENYB[106]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 352.55 0.25 352.65 ;
			LAYER	M2 ;
			RECT	0 352.55 0.25 352.65 ;
			LAYER	M3 ;
			RECT	0 352.55 0.25 352.65 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[106]

	PIN WENYB[107]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 355.43 0.25 355.53 ;
			LAYER	M2 ;
			RECT	0 355.43 0.25 355.53 ;
			LAYER	M3 ;
			RECT	0 355.43 0.25 355.53 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[107]

	PIN WENYB[108]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 358.31 0.25 358.41 ;
			LAYER	M2 ;
			RECT	0 358.31 0.25 358.41 ;
			LAYER	M3 ;
			RECT	0 358.31 0.25 358.41 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[108]

	PIN WENYB[109]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 361.19 0.25 361.29 ;
			LAYER	M2 ;
			RECT	0 361.19 0.25 361.29 ;
			LAYER	M3 ;
			RECT	0 361.19 0.25 361.29 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[109]

	PIN WENYB[10]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.53 0.25 30.63 ;
			LAYER	M2 ;
			RECT	0 30.53 0.25 30.63 ;
			LAYER	M3 ;
			RECT	0 30.53 0.25 30.63 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[10]

	PIN WENYB[110]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 364.07 0.25 364.17 ;
			LAYER	M2 ;
			RECT	0 364.07 0.25 364.17 ;
			LAYER	M3 ;
			RECT	0 364.07 0.25 364.17 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[110]

	PIN WENYB[111]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 366.95 0.25 367.05 ;
			LAYER	M2 ;
			RECT	0 366.95 0.25 367.05 ;
			LAYER	M3 ;
			RECT	0 366.95 0.25 367.05 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[111]

	PIN WENYB[112]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 369.83 0.25 369.93 ;
			LAYER	M2 ;
			RECT	0 369.83 0.25 369.93 ;
			LAYER	M3 ;
			RECT	0 369.83 0.25 369.93 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[112]

	PIN WENYB[113]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 372.71 0.25 372.81 ;
			LAYER	M2 ;
			RECT	0 372.71 0.25 372.81 ;
			LAYER	M3 ;
			RECT	0 372.71 0.25 372.81 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[113]

	PIN WENYB[114]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 375.59 0.25 375.69 ;
			LAYER	M2 ;
			RECT	0 375.59 0.25 375.69 ;
			LAYER	M3 ;
			RECT	0 375.59 0.25 375.69 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[114]

	PIN WENYB[115]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 378.47 0.25 378.57 ;
			LAYER	M2 ;
			RECT	0 378.47 0.25 378.57 ;
			LAYER	M3 ;
			RECT	0 378.47 0.25 378.57 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[115]

	PIN WENYB[116]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 381.35 0.25 381.45 ;
			LAYER	M2 ;
			RECT	0 381.35 0.25 381.45 ;
			LAYER	M3 ;
			RECT	0 381.35 0.25 381.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[116]

	PIN WENYB[117]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 384.23 0.25 384.33 ;
			LAYER	M2 ;
			RECT	0 384.23 0.25 384.33 ;
			LAYER	M3 ;
			RECT	0 384.23 0.25 384.33 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[117]

	PIN WENYB[118]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 387.11 0.25 387.21 ;
			LAYER	M2 ;
			RECT	0 387.11 0.25 387.21 ;
			LAYER	M3 ;
			RECT	0 387.11 0.25 387.21 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[118]

	PIN WENYB[119]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 389.99 0.25 390.09 ;
			LAYER	M2 ;
			RECT	0 389.99 0.25 390.09 ;
			LAYER	M3 ;
			RECT	0 389.99 0.25 390.09 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[119]

	PIN WENYB[11]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.41 0.25 33.51 ;
			LAYER	M2 ;
			RECT	0 33.41 0.25 33.51 ;
			LAYER	M3 ;
			RECT	0 33.41 0.25 33.51 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[11]

	PIN WENYB[120]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 392.87 0.25 392.97 ;
			LAYER	M2 ;
			RECT	0 392.87 0.25 392.97 ;
			LAYER	M3 ;
			RECT	0 392.87 0.25 392.97 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[120]

	PIN WENYB[121]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 395.75 0.25 395.85 ;
			LAYER	M2 ;
			RECT	0 395.75 0.25 395.85 ;
			LAYER	M3 ;
			RECT	0 395.75 0.25 395.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[121]

	PIN WENYB[122]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 398.63 0.25 398.73 ;
			LAYER	M2 ;
			RECT	0 398.63 0.25 398.73 ;
			LAYER	M3 ;
			RECT	0 398.63 0.25 398.73 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[122]

	PIN WENYB[123]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 401.51 0.25 401.61 ;
			LAYER	M2 ;
			RECT	0 401.51 0.25 401.61 ;
			LAYER	M3 ;
			RECT	0 401.51 0.25 401.61 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[123]

	PIN WENYB[124]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 404.39 0.25 404.49 ;
			LAYER	M2 ;
			RECT	0 404.39 0.25 404.49 ;
			LAYER	M3 ;
			RECT	0 404.39 0.25 404.49 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[124]

	PIN WENYB[125]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 407.27 0.25 407.37 ;
			LAYER	M2 ;
			RECT	0 407.27 0.25 407.37 ;
			LAYER	M3 ;
			RECT	0 407.27 0.25 407.37 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[125]

	PIN WENYB[126]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 410.15 0.25 410.25 ;
			LAYER	M2 ;
			RECT	0 410.15 0.25 410.25 ;
			LAYER	M3 ;
			RECT	0 410.15 0.25 410.25 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[126]

	PIN WENYB[127]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 413.03 0.25 413.13 ;
			LAYER	M2 ;
			RECT	0 413.03 0.25 413.13 ;
			LAYER	M3 ;
			RECT	0 413.03 0.25 413.13 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[127]

	PIN WENYB[12]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.29 0.25 36.39 ;
			LAYER	M2 ;
			RECT	0 36.29 0.25 36.39 ;
			LAYER	M3 ;
			RECT	0 36.29 0.25 36.39 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[12]

	PIN WENYB[13]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.17 0.25 39.27 ;
			LAYER	M2 ;
			RECT	0 39.17 0.25 39.27 ;
			LAYER	M3 ;
			RECT	0 39.17 0.25 39.27 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[13]

	PIN WENYB[14]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.05 0.25 42.15 ;
			LAYER	M2 ;
			RECT	0 42.05 0.25 42.15 ;
			LAYER	M3 ;
			RECT	0 42.05 0.25 42.15 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[14]

	PIN WENYB[15]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 44.93 0.25 45.03 ;
			LAYER	M2 ;
			RECT	0 44.93 0.25 45.03 ;
			LAYER	M3 ;
			RECT	0 44.93 0.25 45.03 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[15]

	PIN WENYB[16]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.81 0.25 47.91 ;
			LAYER	M2 ;
			RECT	0 47.81 0.25 47.91 ;
			LAYER	M3 ;
			RECT	0 47.81 0.25 47.91 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[16]

	PIN WENYB[17]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 50.69 0.25 50.79 ;
			LAYER	M2 ;
			RECT	0 50.69 0.25 50.79 ;
			LAYER	M3 ;
			RECT	0 50.69 0.25 50.79 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[17]

	PIN WENYB[18]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 53.57 0.25 53.67 ;
			LAYER	M2 ;
			RECT	0 53.57 0.25 53.67 ;
			LAYER	M3 ;
			RECT	0 53.57 0.25 53.67 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[18]

	PIN WENYB[19]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.45 0.25 56.55 ;
			LAYER	M2 ;
			RECT	0 56.45 0.25 56.55 ;
			LAYER	M3 ;
			RECT	0 56.45 0.25 56.55 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[19]

	PIN WENYB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 4.61 0.25 4.71 ;
			LAYER	M2 ;
			RECT	0 4.61 0.25 4.71 ;
			LAYER	M3 ;
			RECT	0 4.61 0.25 4.71 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[1]

	PIN WENYB[20]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.33 0.25 59.43 ;
			LAYER	M2 ;
			RECT	0 59.33 0.25 59.43 ;
			LAYER	M3 ;
			RECT	0 59.33 0.25 59.43 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[20]

	PIN WENYB[21]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.21 0.25 62.31 ;
			LAYER	M2 ;
			RECT	0 62.21 0.25 62.31 ;
			LAYER	M3 ;
			RECT	0 62.21 0.25 62.31 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[21]

	PIN WENYB[22]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.09 0.25 65.19 ;
			LAYER	M2 ;
			RECT	0 65.09 0.25 65.19 ;
			LAYER	M3 ;
			RECT	0 65.09 0.25 65.19 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[22]

	PIN WENYB[23]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 67.97 0.25 68.07 ;
			LAYER	M2 ;
			RECT	0 67.97 0.25 68.07 ;
			LAYER	M3 ;
			RECT	0 67.97 0.25 68.07 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[23]

	PIN WENYB[24]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 70.85 0.25 70.95 ;
			LAYER	M2 ;
			RECT	0 70.85 0.25 70.95 ;
			LAYER	M3 ;
			RECT	0 70.85 0.25 70.95 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[24]

	PIN WENYB[25]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 73.73 0.25 73.83 ;
			LAYER	M2 ;
			RECT	0 73.73 0.25 73.83 ;
			LAYER	M3 ;
			RECT	0 73.73 0.25 73.83 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[25]

	PIN WENYB[26]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 76.61 0.25 76.71 ;
			LAYER	M2 ;
			RECT	0 76.61 0.25 76.71 ;
			LAYER	M3 ;
			RECT	0 76.61 0.25 76.71 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[26]

	PIN WENYB[27]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.49 0.25 79.59 ;
			LAYER	M2 ;
			RECT	0 79.49 0.25 79.59 ;
			LAYER	M3 ;
			RECT	0 79.49 0.25 79.59 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[27]

	PIN WENYB[28]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.37 0.25 82.47 ;
			LAYER	M2 ;
			RECT	0 82.37 0.25 82.47 ;
			LAYER	M3 ;
			RECT	0 82.37 0.25 82.47 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[28]

	PIN WENYB[29]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 85.25 0.25 85.35 ;
			LAYER	M2 ;
			RECT	0 85.25 0.25 85.35 ;
			LAYER	M3 ;
			RECT	0 85.25 0.25 85.35 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[29]

	PIN WENYB[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.49 0.25 7.59 ;
			LAYER	M2 ;
			RECT	0 7.49 0.25 7.59 ;
			LAYER	M3 ;
			RECT	0 7.49 0.25 7.59 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[2]

	PIN WENYB[30]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 88.13 0.25 88.23 ;
			LAYER	M2 ;
			RECT	0 88.13 0.25 88.23 ;
			LAYER	M3 ;
			RECT	0 88.13 0.25 88.23 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[30]

	PIN WENYB[31]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 91.01 0.25 91.11 ;
			LAYER	M2 ;
			RECT	0 91.01 0.25 91.11 ;
			LAYER	M3 ;
			RECT	0 91.01 0.25 91.11 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[31]

	PIN WENYB[32]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 93.89 0.25 93.99 ;
			LAYER	M2 ;
			RECT	0 93.89 0.25 93.99 ;
			LAYER	M3 ;
			RECT	0 93.89 0.25 93.99 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[32]

	PIN WENYB[33]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 96.77 0.25 96.87 ;
			LAYER	M2 ;
			RECT	0 96.77 0.25 96.87 ;
			LAYER	M3 ;
			RECT	0 96.77 0.25 96.87 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[33]

	PIN WENYB[34]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 99.65 0.25 99.75 ;
			LAYER	M2 ;
			RECT	0 99.65 0.25 99.75 ;
			LAYER	M3 ;
			RECT	0 99.65 0.25 99.75 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[34]

	PIN WENYB[35]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 102.53 0.25 102.63 ;
			LAYER	M2 ;
			RECT	0 102.53 0.25 102.63 ;
			LAYER	M3 ;
			RECT	0 102.53 0.25 102.63 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[35]

	PIN WENYB[36]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 105.41 0.25 105.51 ;
			LAYER	M2 ;
			RECT	0 105.41 0.25 105.51 ;
			LAYER	M3 ;
			RECT	0 105.41 0.25 105.51 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[36]

	PIN WENYB[37]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 108.29 0.25 108.39 ;
			LAYER	M2 ;
			RECT	0 108.29 0.25 108.39 ;
			LAYER	M3 ;
			RECT	0 108.29 0.25 108.39 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[37]

	PIN WENYB[38]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 111.17 0.25 111.27 ;
			LAYER	M2 ;
			RECT	0 111.17 0.25 111.27 ;
			LAYER	M3 ;
			RECT	0 111.17 0.25 111.27 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[38]

	PIN WENYB[39]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 114.05 0.25 114.15 ;
			LAYER	M2 ;
			RECT	0 114.05 0.25 114.15 ;
			LAYER	M3 ;
			RECT	0 114.05 0.25 114.15 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[39]

	PIN WENYB[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.37 0.25 10.47 ;
			LAYER	M2 ;
			RECT	0 10.37 0.25 10.47 ;
			LAYER	M3 ;
			RECT	0 10.37 0.25 10.47 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[3]

	PIN WENYB[40]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 116.93 0.25 117.03 ;
			LAYER	M2 ;
			RECT	0 116.93 0.25 117.03 ;
			LAYER	M3 ;
			RECT	0 116.93 0.25 117.03 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[40]

	PIN WENYB[41]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 119.81 0.25 119.91 ;
			LAYER	M2 ;
			RECT	0 119.81 0.25 119.91 ;
			LAYER	M3 ;
			RECT	0 119.81 0.25 119.91 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[41]

	PIN WENYB[42]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 122.69 0.25 122.79 ;
			LAYER	M2 ;
			RECT	0 122.69 0.25 122.79 ;
			LAYER	M3 ;
			RECT	0 122.69 0.25 122.79 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[42]

	PIN WENYB[43]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 125.57 0.25 125.67 ;
			LAYER	M2 ;
			RECT	0 125.57 0.25 125.67 ;
			LAYER	M3 ;
			RECT	0 125.57 0.25 125.67 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[43]

	PIN WENYB[44]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 128.45 0.25 128.55 ;
			LAYER	M2 ;
			RECT	0 128.45 0.25 128.55 ;
			LAYER	M3 ;
			RECT	0 128.45 0.25 128.55 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[44]

	PIN WENYB[45]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 131.33 0.25 131.43 ;
			LAYER	M2 ;
			RECT	0 131.33 0.25 131.43 ;
			LAYER	M3 ;
			RECT	0 131.33 0.25 131.43 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[45]

	PIN WENYB[46]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 134.21 0.25 134.31 ;
			LAYER	M2 ;
			RECT	0 134.21 0.25 134.31 ;
			LAYER	M3 ;
			RECT	0 134.21 0.25 134.31 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[46]

	PIN WENYB[47]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 137.09 0.25 137.19 ;
			LAYER	M2 ;
			RECT	0 137.09 0.25 137.19 ;
			LAYER	M3 ;
			RECT	0 137.09 0.25 137.19 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[47]

	PIN WENYB[48]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 139.97 0.25 140.07 ;
			LAYER	M2 ;
			RECT	0 139.97 0.25 140.07 ;
			LAYER	M3 ;
			RECT	0 139.97 0.25 140.07 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[48]

	PIN WENYB[49]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 142.85 0.25 142.95 ;
			LAYER	M2 ;
			RECT	0 142.85 0.25 142.95 ;
			LAYER	M3 ;
			RECT	0 142.85 0.25 142.95 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[49]

	PIN WENYB[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.25 0.25 13.35 ;
			LAYER	M2 ;
			RECT	0 13.25 0.25 13.35 ;
			LAYER	M3 ;
			RECT	0 13.25 0.25 13.35 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[4]

	PIN WENYB[50]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 145.73 0.25 145.83 ;
			LAYER	M2 ;
			RECT	0 145.73 0.25 145.83 ;
			LAYER	M3 ;
			RECT	0 145.73 0.25 145.83 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[50]

	PIN WENYB[51]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 148.61 0.25 148.71 ;
			LAYER	M2 ;
			RECT	0 148.61 0.25 148.71 ;
			LAYER	M3 ;
			RECT	0 148.61 0.25 148.71 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[51]

	PIN WENYB[52]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 151.49 0.25 151.59 ;
			LAYER	M2 ;
			RECT	0 151.49 0.25 151.59 ;
			LAYER	M3 ;
			RECT	0 151.49 0.25 151.59 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[52]

	PIN WENYB[53]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 154.37 0.25 154.47 ;
			LAYER	M2 ;
			RECT	0 154.37 0.25 154.47 ;
			LAYER	M3 ;
			RECT	0 154.37 0.25 154.47 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[53]

	PIN WENYB[54]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 157.25 0.25 157.35 ;
			LAYER	M2 ;
			RECT	0 157.25 0.25 157.35 ;
			LAYER	M3 ;
			RECT	0 157.25 0.25 157.35 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[54]

	PIN WENYB[55]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 160.13 0.25 160.23 ;
			LAYER	M2 ;
			RECT	0 160.13 0.25 160.23 ;
			LAYER	M3 ;
			RECT	0 160.13 0.25 160.23 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[55]

	PIN WENYB[56]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 163.01 0.25 163.11 ;
			LAYER	M2 ;
			RECT	0 163.01 0.25 163.11 ;
			LAYER	M3 ;
			RECT	0 163.01 0.25 163.11 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[56]

	PIN WENYB[57]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 165.89 0.25 165.99 ;
			LAYER	M2 ;
			RECT	0 165.89 0.25 165.99 ;
			LAYER	M3 ;
			RECT	0 165.89 0.25 165.99 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[57]

	PIN WENYB[58]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 168.77 0.25 168.87 ;
			LAYER	M2 ;
			RECT	0 168.77 0.25 168.87 ;
			LAYER	M3 ;
			RECT	0 168.77 0.25 168.87 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[58]

	PIN WENYB[59]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 171.65 0.25 171.75 ;
			LAYER	M2 ;
			RECT	0 171.65 0.25 171.75 ;
			LAYER	M3 ;
			RECT	0 171.65 0.25 171.75 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[59]

	PIN WENYB[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.13 0.25 16.23 ;
			LAYER	M2 ;
			RECT	0 16.13 0.25 16.23 ;
			LAYER	M3 ;
			RECT	0 16.13 0.25 16.23 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[5]

	PIN WENYB[60]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 174.53 0.25 174.63 ;
			LAYER	M2 ;
			RECT	0 174.53 0.25 174.63 ;
			LAYER	M3 ;
			RECT	0 174.53 0.25 174.63 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[60]

	PIN WENYB[61]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 177.41 0.25 177.51 ;
			LAYER	M2 ;
			RECT	0 177.41 0.25 177.51 ;
			LAYER	M3 ;
			RECT	0 177.41 0.25 177.51 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[61]

	PIN WENYB[62]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 180.29 0.25 180.39 ;
			LAYER	M2 ;
			RECT	0 180.29 0.25 180.39 ;
			LAYER	M3 ;
			RECT	0 180.29 0.25 180.39 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[62]

	PIN WENYB[63]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 183.17 0.25 183.27 ;
			LAYER	M2 ;
			RECT	0 183.17 0.25 183.27 ;
			LAYER	M3 ;
			RECT	0 183.17 0.25 183.27 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[63]

	PIN WENYB[64]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 231.59 0.25 231.69 ;
			LAYER	M2 ;
			RECT	0 231.59 0.25 231.69 ;
			LAYER	M3 ;
			RECT	0 231.59 0.25 231.69 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[64]

	PIN WENYB[65]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 234.47 0.25 234.57 ;
			LAYER	M2 ;
			RECT	0 234.47 0.25 234.57 ;
			LAYER	M3 ;
			RECT	0 234.47 0.25 234.57 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[65]

	PIN WENYB[66]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 237.35 0.25 237.45 ;
			LAYER	M2 ;
			RECT	0 237.35 0.25 237.45 ;
			LAYER	M3 ;
			RECT	0 237.35 0.25 237.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[66]

	PIN WENYB[67]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 240.23 0.25 240.33 ;
			LAYER	M2 ;
			RECT	0 240.23 0.25 240.33 ;
			LAYER	M3 ;
			RECT	0 240.23 0.25 240.33 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[67]

	PIN WENYB[68]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 243.11 0.25 243.21 ;
			LAYER	M2 ;
			RECT	0 243.11 0.25 243.21 ;
			LAYER	M3 ;
			RECT	0 243.11 0.25 243.21 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[68]

	PIN WENYB[69]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 245.99 0.25 246.09 ;
			LAYER	M2 ;
			RECT	0 245.99 0.25 246.09 ;
			LAYER	M3 ;
			RECT	0 245.99 0.25 246.09 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[69]

	PIN WENYB[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.01 0.25 19.11 ;
			LAYER	M2 ;
			RECT	0 19.01 0.25 19.11 ;
			LAYER	M3 ;
			RECT	0 19.01 0.25 19.11 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[6]

	PIN WENYB[70]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 248.87 0.25 248.97 ;
			LAYER	M2 ;
			RECT	0 248.87 0.25 248.97 ;
			LAYER	M3 ;
			RECT	0 248.87 0.25 248.97 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[70]

	PIN WENYB[71]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 251.75 0.25 251.85 ;
			LAYER	M2 ;
			RECT	0 251.75 0.25 251.85 ;
			LAYER	M3 ;
			RECT	0 251.75 0.25 251.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[71]

	PIN WENYB[72]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 254.63 0.25 254.73 ;
			LAYER	M2 ;
			RECT	0 254.63 0.25 254.73 ;
			LAYER	M3 ;
			RECT	0 254.63 0.25 254.73 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[72]

	PIN WENYB[73]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 257.51 0.25 257.61 ;
			LAYER	M2 ;
			RECT	0 257.51 0.25 257.61 ;
			LAYER	M3 ;
			RECT	0 257.51 0.25 257.61 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[73]

	PIN WENYB[74]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 260.39 0.25 260.49 ;
			LAYER	M2 ;
			RECT	0 260.39 0.25 260.49 ;
			LAYER	M3 ;
			RECT	0 260.39 0.25 260.49 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[74]

	PIN WENYB[75]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 263.27 0.25 263.37 ;
			LAYER	M2 ;
			RECT	0 263.27 0.25 263.37 ;
			LAYER	M3 ;
			RECT	0 263.27 0.25 263.37 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[75]

	PIN WENYB[76]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 266.15 0.25 266.25 ;
			LAYER	M2 ;
			RECT	0 266.15 0.25 266.25 ;
			LAYER	M3 ;
			RECT	0 266.15 0.25 266.25 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[76]

	PIN WENYB[77]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 269.03 0.25 269.13 ;
			LAYER	M2 ;
			RECT	0 269.03 0.25 269.13 ;
			LAYER	M3 ;
			RECT	0 269.03 0.25 269.13 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[77]

	PIN WENYB[78]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 271.91 0.25 272.01 ;
			LAYER	M2 ;
			RECT	0 271.91 0.25 272.01 ;
			LAYER	M3 ;
			RECT	0 271.91 0.25 272.01 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[78]

	PIN WENYB[79]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 274.79 0.25 274.89 ;
			LAYER	M2 ;
			RECT	0 274.79 0.25 274.89 ;
			LAYER	M3 ;
			RECT	0 274.79 0.25 274.89 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[79]

	PIN WENYB[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 21.89 0.25 21.99 ;
			LAYER	M2 ;
			RECT	0 21.89 0.25 21.99 ;
			LAYER	M3 ;
			RECT	0 21.89 0.25 21.99 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[7]

	PIN WENYB[80]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 277.67 0.25 277.77 ;
			LAYER	M2 ;
			RECT	0 277.67 0.25 277.77 ;
			LAYER	M3 ;
			RECT	0 277.67 0.25 277.77 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[80]

	PIN WENYB[81]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 280.55 0.25 280.65 ;
			LAYER	M2 ;
			RECT	0 280.55 0.25 280.65 ;
			LAYER	M3 ;
			RECT	0 280.55 0.25 280.65 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[81]

	PIN WENYB[82]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 283.43 0.25 283.53 ;
			LAYER	M2 ;
			RECT	0 283.43 0.25 283.53 ;
			LAYER	M3 ;
			RECT	0 283.43 0.25 283.53 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[82]

	PIN WENYB[83]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 286.31 0.25 286.41 ;
			LAYER	M2 ;
			RECT	0 286.31 0.25 286.41 ;
			LAYER	M3 ;
			RECT	0 286.31 0.25 286.41 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[83]

	PIN WENYB[84]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 289.19 0.25 289.29 ;
			LAYER	M2 ;
			RECT	0 289.19 0.25 289.29 ;
			LAYER	M3 ;
			RECT	0 289.19 0.25 289.29 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[84]

	PIN WENYB[85]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 292.07 0.25 292.17 ;
			LAYER	M2 ;
			RECT	0 292.07 0.25 292.17 ;
			LAYER	M3 ;
			RECT	0 292.07 0.25 292.17 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[85]

	PIN WENYB[86]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 294.95 0.25 295.05 ;
			LAYER	M2 ;
			RECT	0 294.95 0.25 295.05 ;
			LAYER	M3 ;
			RECT	0 294.95 0.25 295.05 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[86]

	PIN WENYB[87]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 297.83 0.25 297.93 ;
			LAYER	M2 ;
			RECT	0 297.83 0.25 297.93 ;
			LAYER	M3 ;
			RECT	0 297.83 0.25 297.93 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[87]

	PIN WENYB[88]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 300.71 0.25 300.81 ;
			LAYER	M2 ;
			RECT	0 300.71 0.25 300.81 ;
			LAYER	M3 ;
			RECT	0 300.71 0.25 300.81 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[88]

	PIN WENYB[89]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 303.59 0.25 303.69 ;
			LAYER	M2 ;
			RECT	0 303.59 0.25 303.69 ;
			LAYER	M3 ;
			RECT	0 303.59 0.25 303.69 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[89]

	PIN WENYB[8]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 24.77 0.25 24.87 ;
			LAYER	M2 ;
			RECT	0 24.77 0.25 24.87 ;
			LAYER	M3 ;
			RECT	0 24.77 0.25 24.87 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[8]

	PIN WENYB[90]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 306.47 0.25 306.57 ;
			LAYER	M2 ;
			RECT	0 306.47 0.25 306.57 ;
			LAYER	M3 ;
			RECT	0 306.47 0.25 306.57 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[90]

	PIN WENYB[91]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 309.35 0.25 309.45 ;
			LAYER	M2 ;
			RECT	0 309.35 0.25 309.45 ;
			LAYER	M3 ;
			RECT	0 309.35 0.25 309.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[91]

	PIN WENYB[92]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 312.23 0.25 312.33 ;
			LAYER	M2 ;
			RECT	0 312.23 0.25 312.33 ;
			LAYER	M3 ;
			RECT	0 312.23 0.25 312.33 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[92]

	PIN WENYB[93]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 315.11 0.25 315.21 ;
			LAYER	M2 ;
			RECT	0 315.11 0.25 315.21 ;
			LAYER	M3 ;
			RECT	0 315.11 0.25 315.21 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[93]

	PIN WENYB[94]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 317.99 0.25 318.09 ;
			LAYER	M2 ;
			RECT	0 317.99 0.25 318.09 ;
			LAYER	M3 ;
			RECT	0 317.99 0.25 318.09 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[94]

	PIN WENYB[95]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 320.87 0.25 320.97 ;
			LAYER	M2 ;
			RECT	0 320.87 0.25 320.97 ;
			LAYER	M3 ;
			RECT	0 320.87 0.25 320.97 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[95]

	PIN WENYB[96]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 323.75 0.25 323.85 ;
			LAYER	M2 ;
			RECT	0 323.75 0.25 323.85 ;
			LAYER	M3 ;
			RECT	0 323.75 0.25 323.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[96]

	PIN WENYB[97]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 326.63 0.25 326.73 ;
			LAYER	M2 ;
			RECT	0 326.63 0.25 326.73 ;
			LAYER	M3 ;
			RECT	0 326.63 0.25 326.73 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[97]

	PIN WENYB[98]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 329.51 0.25 329.61 ;
			LAYER	M2 ;
			RECT	0 329.51 0.25 329.61 ;
			LAYER	M3 ;
			RECT	0 329.51 0.25 329.61 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[98]

	PIN WENYB[99]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 332.39 0.25 332.49 ;
			LAYER	M2 ;
			RECT	0 332.39 0.25 332.49 ;
			LAYER	M3 ;
			RECT	0 332.39 0.25 332.49 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[99]

	PIN WENYB[9]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 27.65 0.25 27.75 ;
			LAYER	M2 ;
			RECT	0 27.65 0.25 27.75 ;
			LAYER	M3 ;
			RECT	0 27.65 0.25 27.75 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[9]

	OBS
		LAYER	M1 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 20.845 414.51 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 2.655 0.32 3.16 ;
		RECT	0 3.46 0.32 4.245 ;
		RECT	0 5.535 0.32 6.04 ;
		RECT	0 6.34 0.32 7.125 ;
		RECT	0 8.415 0.32 8.92 ;
		RECT	0 9.22 0.32 10.005 ;
		RECT	0 11.295 0.32 11.8 ;
		RECT	0 12.1 0.32 12.885 ;
		RECT	0 14.175 0.32 14.68 ;
		RECT	0 14.98 0.32 15.765 ;
		RECT	0 17.055 0.32 17.56 ;
		RECT	0 17.86 0.32 18.645 ;
		RECT	0 19.935 0.32 20.44 ;
		RECT	0 20.74 0.32 21.525 ;
		RECT	0 22.815 0.32 23.32 ;
		RECT	0 23.62 0.32 24.405 ;
		RECT	0 25.695 0.32 26.2 ;
		RECT	0 26.5 0.32 27.285 ;
		RECT	0 28.575 0.32 29.08 ;
		RECT	0 29.38 0.32 30.165 ;
		RECT	0 31.455 0.32 31.96 ;
		RECT	0 32.26 0.32 33.045 ;
		RECT	0 34.335 0.32 34.84 ;
		RECT	0 35.14 0.32 35.925 ;
		RECT	0 37.215 0.32 37.72 ;
		RECT	0 38.02 0.32 38.805 ;
		RECT	0 40.095 0.32 40.6 ;
		RECT	0 40.9 0.32 41.685 ;
		RECT	0 42.975 0.32 43.48 ;
		RECT	0 43.78 0.32 44.565 ;
		RECT	0 45.855 0.32 46.36 ;
		RECT	0 46.66 0.32 47.445 ;
		RECT	0 48.735 0.32 49.24 ;
		RECT	0 49.54 0.32 50.325 ;
		RECT	0 51.615 0.32 52.12 ;
		RECT	0 52.42 0.32 53.205 ;
		RECT	0 54.495 0.32 55 ;
		RECT	0 55.3 0.32 56.085 ;
		RECT	0 57.375 0.32 57.88 ;
		RECT	0 58.18 0.32 58.965 ;
		RECT	0 60.255 0.32 60.76 ;
		RECT	0 61.06 0.32 61.845 ;
		RECT	0 63.135 0.32 63.64 ;
		RECT	0 63.94 0.32 64.725 ;
		RECT	0 66.015 0.32 66.52 ;
		RECT	0 66.82 0.32 67.605 ;
		RECT	0 68.895 0.32 69.4 ;
		RECT	0 69.7 0.32 70.485 ;
		RECT	0 71.775 0.32 72.28 ;
		RECT	0 72.58 0.32 73.365 ;
		RECT	0 74.655 0.32 75.16 ;
		RECT	0 75.46 0.32 76.245 ;
		RECT	0 77.535 0.32 78.04 ;
		RECT	0 78.34 0.32 79.125 ;
		RECT	0 80.415 0.32 80.92 ;
		RECT	0 81.22 0.32 82.005 ;
		RECT	0 83.295 0.32 83.8 ;
		RECT	0 84.1 0.32 84.885 ;
		RECT	0 86.175 0.32 86.68 ;
		RECT	0 86.98 0.32 87.765 ;
		RECT	0 89.055 0.32 89.56 ;
		RECT	0 89.86 0.32 90.645 ;
		RECT	0 91.935 0.32 92.44 ;
		RECT	0 92.74 0.32 93.525 ;
		RECT	0 94.815 0.32 95.32 ;
		RECT	0 95.62 0.32 96.405 ;
		RECT	0 97.695 0.32 98.2 ;
		RECT	0 98.5 0.32 99.285 ;
		RECT	0 100.575 0.32 101.08 ;
		RECT	0 101.38 0.32 102.165 ;
		RECT	0 103.455 0.32 103.96 ;
		RECT	0 104.26 0.32 105.045 ;
		RECT	0 106.335 0.32 106.84 ;
		RECT	0 107.14 0.32 107.925 ;
		RECT	0 109.215 0.32 109.72 ;
		RECT	0 110.02 0.32 110.805 ;
		RECT	0 112.095 0.32 112.6 ;
		RECT	0 112.9 0.32 113.685 ;
		RECT	0 114.975 0.32 115.48 ;
		RECT	0 115.78 0.32 116.565 ;
		RECT	0 117.855 0.32 118.36 ;
		RECT	0 118.66 0.32 119.445 ;
		RECT	0 120.735 0.32 121.24 ;
		RECT	0 121.54 0.32 122.325 ;
		RECT	0 123.615 0.32 124.12 ;
		RECT	0 124.42 0.32 125.205 ;
		RECT	0 126.495 0.32 127 ;
		RECT	0 127.3 0.32 128.085 ;
		RECT	0 129.375 0.32 129.88 ;
		RECT	0 130.18 0.32 130.965 ;
		RECT	0 132.255 0.32 132.76 ;
		RECT	0 133.06 0.32 133.845 ;
		RECT	0 135.135 0.32 135.64 ;
		RECT	0 135.94 0.32 136.725 ;
		RECT	0 138.015 0.32 138.52 ;
		RECT	0 138.82 0.32 139.605 ;
		RECT	0 140.895 0.32 141.4 ;
		RECT	0 141.7 0.32 142.485 ;
		RECT	0 143.775 0.32 144.28 ;
		RECT	0 144.58 0.32 145.365 ;
		RECT	0 146.655 0.32 147.16 ;
		RECT	0 147.46 0.32 148.245 ;
		RECT	0 149.535 0.32 150.04 ;
		RECT	0 150.34 0.32 151.125 ;
		RECT	0 152.415 0.32 152.92 ;
		RECT	0 153.22 0.32 154.005 ;
		RECT	0 155.295 0.32 155.8 ;
		RECT	0 156.1 0.32 156.885 ;
		RECT	0 158.175 0.32 158.68 ;
		RECT	0 158.98 0.32 159.765 ;
		RECT	0 161.055 0.32 161.56 ;
		RECT	0 161.86 0.32 162.645 ;
		RECT	0 163.935 0.32 164.44 ;
		RECT	0 164.74 0.32 165.525 ;
		RECT	0 166.815 0.32 167.32 ;
		RECT	0 167.62 0.32 168.405 ;
		RECT	0 169.695 0.32 170.2 ;
		RECT	0 170.5 0.32 171.285 ;
		RECT	0 172.575 0.32 173.08 ;
		RECT	0 173.38 0.32 174.165 ;
		RECT	0 175.455 0.32 175.96 ;
		RECT	0 176.26 0.32 177.045 ;
		RECT	0 178.335 0.32 178.84 ;
		RECT	0 179.14 0.32 179.925 ;
		RECT	0 181.215 0.32 181.72 ;
		RECT	0 182.02 0.32 182.805 ;
		RECT	0 184.095 0.32 184.6 ;
		RECT	0 184.9 0.32 187 ;
		RECT	0 187.3 0.32 187.35 ;
		RECT	0 187.65 0.32 188.01 ;
		RECT	0 188.71 0.32 190.35 ;
		RECT	0 190.955 0.32 191.17 ;
		RECT	0 191.47 0.32 191.575 ;
		RECT	0 191.875 0.32 193.685 ;
		RECT	0 193.985 0.32 194.2 ;
		RECT	0 194.5 0.32 194.605 ;
		RECT	0 194.905 0.32 196.745 ;
		RECT	0 197.045 0.32 197.23 ;
		RECT	0 197.53 0.32 197.635 ;
		RECT	0 197.935 0.32 198.03 ;
		RECT	0 198.33 0.32 198.4 ;
		RECT	0 198.7 0.32 198.775 ;
		RECT	0 199.075 0.32 199.26 ;
		RECT	0 199.97 0.32 201.405 ;
		RECT	0 202.105 0.32 202.29 ;
		RECT	0 202.875 0.32 205.8 ;
		RECT	0 206.5 0.32 206.97 ;
		RECT	0 207.27 0.32 208.635 ;
		RECT	0 208.935 0.32 212.725 ;
		RECT	0 213.26 0.32 213.45 ;
		RECT	0 213.75 0.32 213.825 ;
		RECT	0 214.125 0.32 214.205 ;
		RECT	0 214.505 0.32 215.205 ;
		RECT	0 215.505 0.32 215.995 ;
		RECT	0 216.295 0.32 216.48 ;
		RECT	0 216.78 0.32 216.885 ;
		RECT	0 217.185 0.32 217.65 ;
		RECT	0 217.95 0.32 218.025 ;
		RECT	0 218.325 0.32 218.48 ;
		RECT	0 218.98 0.32 220.225 ;
		RECT	0 220.525 0.32 220.65 ;
		RECT	0 221.16 0.32 221.54 ;
		RECT	0 221.84 0.32 223.68 ;
		RECT	0 223.98 0.32 224.085 ;
		RECT	0 224.385 0.32 224.57 ;
		RECT	0 225.125 0.32 225.6 ;
		RECT	0 225.9 0.32 228.21 ;
		RECT	0 228.51 0.32 228.605 ;
		RECT	0 228.905 0.32 229.15 ;
		RECT	0 229.45 0.32 229.96 ;
		RECT	0 230.26 0.32 230.765 ;
		RECT	0 232.055 0.32 232.84 ;
		RECT	0 233.14 0.32 233.645 ;
		RECT	0 234.935 0.32 235.72 ;
		RECT	0 236.02 0.32 236.525 ;
		RECT	0 237.815 0.32 238.6 ;
		RECT	0 238.9 0.32 239.405 ;
		RECT	0 240.695 0.32 241.48 ;
		RECT	0 241.78 0.32 242.285 ;
		RECT	0 243.575 0.32 244.36 ;
		RECT	0 244.66 0.32 245.165 ;
		RECT	0 246.455 0.32 247.24 ;
		RECT	0 247.54 0.32 248.045 ;
		RECT	0 249.335 0.32 250.12 ;
		RECT	0 250.42 0.32 250.925 ;
		RECT	0 252.215 0.32 253 ;
		RECT	0 253.3 0.32 253.805 ;
		RECT	0 255.095 0.32 255.88 ;
		RECT	0 256.18 0.32 256.685 ;
		RECT	0 257.975 0.32 258.76 ;
		RECT	0 259.06 0.32 259.565 ;
		RECT	0 260.855 0.32 261.64 ;
		RECT	0 261.94 0.32 262.445 ;
		RECT	0 263.735 0.32 264.52 ;
		RECT	0 264.82 0.32 265.325 ;
		RECT	0 266.615 0.32 267.4 ;
		RECT	0 267.7 0.32 268.205 ;
		RECT	0 269.495 0.32 270.28 ;
		RECT	0 270.58 0.32 271.085 ;
		RECT	0 272.375 0.32 273.16 ;
		RECT	0 273.46 0.32 273.965 ;
		RECT	0 275.255 0.32 276.04 ;
		RECT	0 276.34 0.32 276.845 ;
		RECT	0 278.135 0.32 278.92 ;
		RECT	0 279.22 0.32 279.725 ;
		RECT	0 281.015 0.32 281.8 ;
		RECT	0 282.1 0.32 282.605 ;
		RECT	0 283.895 0.32 284.68 ;
		RECT	0 284.98 0.32 285.485 ;
		RECT	0 286.775 0.32 287.56 ;
		RECT	0 287.86 0.32 288.365 ;
		RECT	0 289.655 0.32 290.44 ;
		RECT	0 290.74 0.32 291.245 ;
		RECT	0 292.535 0.32 293.32 ;
		RECT	0 293.62 0.32 294.125 ;
		RECT	0 295.415 0.32 296.2 ;
		RECT	0 296.5 0.32 297.005 ;
		RECT	0 298.295 0.32 299.08 ;
		RECT	0 299.38 0.32 299.885 ;
		RECT	0 301.175 0.32 301.96 ;
		RECT	0 302.26 0.32 302.765 ;
		RECT	0 304.055 0.32 304.84 ;
		RECT	0 305.14 0.32 305.645 ;
		RECT	0 306.935 0.32 307.72 ;
		RECT	0 308.02 0.32 308.525 ;
		RECT	0 309.815 0.32 310.6 ;
		RECT	0 310.9 0.32 311.405 ;
		RECT	0 312.695 0.32 313.48 ;
		RECT	0 313.78 0.32 314.285 ;
		RECT	0 315.575 0.32 316.36 ;
		RECT	0 316.66 0.32 317.165 ;
		RECT	0 318.455 0.32 319.24 ;
		RECT	0 319.54 0.32 320.045 ;
		RECT	0 321.335 0.32 322.12 ;
		RECT	0 322.42 0.32 322.925 ;
		RECT	0 324.215 0.32 325 ;
		RECT	0 325.3 0.32 325.805 ;
		RECT	0 327.095 0.32 327.88 ;
		RECT	0 328.18 0.32 328.685 ;
		RECT	0 329.975 0.32 330.76 ;
		RECT	0 331.06 0.32 331.565 ;
		RECT	0 332.855 0.32 333.64 ;
		RECT	0 333.94 0.32 334.445 ;
		RECT	0 335.735 0.32 336.52 ;
		RECT	0 336.82 0.32 337.325 ;
		RECT	0 338.615 0.32 339.4 ;
		RECT	0 339.7 0.32 340.205 ;
		RECT	0 341.495 0.32 342.28 ;
		RECT	0 342.58 0.32 343.085 ;
		RECT	0 344.375 0.32 345.16 ;
		RECT	0 345.46 0.32 345.965 ;
		RECT	0 347.255 0.32 348.04 ;
		RECT	0 348.34 0.32 348.845 ;
		RECT	0 350.135 0.32 350.92 ;
		RECT	0 351.22 0.32 351.725 ;
		RECT	0 353.015 0.32 353.8 ;
		RECT	0 354.1 0.32 354.605 ;
		RECT	0 355.895 0.32 356.68 ;
		RECT	0 356.98 0.32 357.485 ;
		RECT	0 358.775 0.32 359.56 ;
		RECT	0 359.86 0.32 360.365 ;
		RECT	0 361.655 0.32 362.44 ;
		RECT	0 362.74 0.32 363.245 ;
		RECT	0 364.535 0.32 365.32 ;
		RECT	0 365.62 0.32 366.125 ;
		RECT	0 367.415 0.32 368.2 ;
		RECT	0 368.5 0.32 369.005 ;
		RECT	0 370.295 0.32 371.08 ;
		RECT	0 371.38 0.32 371.885 ;
		RECT	0 373.175 0.32 373.96 ;
		RECT	0 374.26 0.32 374.765 ;
		RECT	0 376.055 0.32 376.84 ;
		RECT	0 377.14 0.32 377.645 ;
		RECT	0 378.935 0.32 379.72 ;
		RECT	0 380.02 0.32 380.525 ;
		RECT	0 381.815 0.32 382.6 ;
		RECT	0 382.9 0.32 383.405 ;
		RECT	0 384.695 0.32 385.48 ;
		RECT	0 385.78 0.32 386.285 ;
		RECT	0 387.575 0.32 388.36 ;
		RECT	0 388.66 0.32 389.165 ;
		RECT	0 390.455 0.32 391.24 ;
		RECT	0 391.54 0.32 392.045 ;
		RECT	0 393.335 0.32 394.12 ;
		RECT	0 394.42 0.32 394.925 ;
		RECT	0 396.215 0.32 397 ;
		RECT	0 397.3 0.32 397.805 ;
		RECT	0 399.095 0.32 399.88 ;
		RECT	0 400.18 0.32 400.685 ;
		RECT	0 401.975 0.32 402.76 ;
		RECT	0 403.06 0.32 403.565 ;
		RECT	0 404.855 0.32 405.64 ;
		RECT	0 405.94 0.32 406.445 ;
		RECT	0 407.735 0.32 408.52 ;
		RECT	0 408.82 0.32 409.325 ;
		RECT	0 410.615 0.32 411.4 ;
		RECT	0 411.7 0.32 412.205 ;
		RECT	0 413.495 0.32 414.3 ;
		RECT	20.845 0 21.165 414.86 ;
		RECT	0.32 0 20.845 0.35 ;
		RECT	0.32 414.51 20.845 414.86 ;
		LAYER	M2 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 20.845 414.51 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 2.655 0.32 3.16 ;
		RECT	0 3.46 0.32 4.245 ;
		RECT	0 5.535 0.32 6.04 ;
		RECT	0 6.34 0.32 7.125 ;
		RECT	0 8.415 0.32 8.92 ;
		RECT	0 9.22 0.32 10.005 ;
		RECT	0 11.295 0.32 11.8 ;
		RECT	0 12.1 0.32 12.885 ;
		RECT	0 14.175 0.32 14.68 ;
		RECT	0 14.98 0.32 15.765 ;
		RECT	0 17.055 0.32 17.56 ;
		RECT	0 17.86 0.32 18.645 ;
		RECT	0 19.935 0.32 20.44 ;
		RECT	0 20.74 0.32 21.525 ;
		RECT	0 22.815 0.32 23.32 ;
		RECT	0 23.62 0.32 24.405 ;
		RECT	0 25.695 0.32 26.2 ;
		RECT	0 26.5 0.32 27.285 ;
		RECT	0 28.575 0.32 29.08 ;
		RECT	0 29.38 0.32 30.165 ;
		RECT	0 31.455 0.32 31.96 ;
		RECT	0 32.26 0.32 33.045 ;
		RECT	0 34.335 0.32 34.84 ;
		RECT	0 35.14 0.32 35.925 ;
		RECT	0 37.215 0.32 37.72 ;
		RECT	0 38.02 0.32 38.805 ;
		RECT	0 40.095 0.32 40.6 ;
		RECT	0 40.9 0.32 41.685 ;
		RECT	0 42.975 0.32 43.48 ;
		RECT	0 43.78 0.32 44.565 ;
		RECT	0 45.855 0.32 46.36 ;
		RECT	0 46.66 0.32 47.445 ;
		RECT	0 48.735 0.32 49.24 ;
		RECT	0 49.54 0.32 50.325 ;
		RECT	0 51.615 0.32 52.12 ;
		RECT	0 52.42 0.32 53.205 ;
		RECT	0 54.495 0.32 55 ;
		RECT	0 55.3 0.32 56.085 ;
		RECT	0 57.375 0.32 57.88 ;
		RECT	0 58.18 0.32 58.965 ;
		RECT	0 60.255 0.32 60.76 ;
		RECT	0 61.06 0.32 61.845 ;
		RECT	0 63.135 0.32 63.64 ;
		RECT	0 63.94 0.32 64.725 ;
		RECT	0 66.015 0.32 66.52 ;
		RECT	0 66.82 0.32 67.605 ;
		RECT	0 68.895 0.32 69.4 ;
		RECT	0 69.7 0.32 70.485 ;
		RECT	0 71.775 0.32 72.28 ;
		RECT	0 72.58 0.32 73.365 ;
		RECT	0 74.655 0.32 75.16 ;
		RECT	0 75.46 0.32 76.245 ;
		RECT	0 77.535 0.32 78.04 ;
		RECT	0 78.34 0.32 79.125 ;
		RECT	0 80.415 0.32 80.92 ;
		RECT	0 81.22 0.32 82.005 ;
		RECT	0 83.295 0.32 83.8 ;
		RECT	0 84.1 0.32 84.885 ;
		RECT	0 86.175 0.32 86.68 ;
		RECT	0 86.98 0.32 87.765 ;
		RECT	0 89.055 0.32 89.56 ;
		RECT	0 89.86 0.32 90.645 ;
		RECT	0 91.935 0.32 92.44 ;
		RECT	0 92.74 0.32 93.525 ;
		RECT	0 94.815 0.32 95.32 ;
		RECT	0 95.62 0.32 96.405 ;
		RECT	0 97.695 0.32 98.2 ;
		RECT	0 98.5 0.32 99.285 ;
		RECT	0 100.575 0.32 101.08 ;
		RECT	0 101.38 0.32 102.165 ;
		RECT	0 103.455 0.32 103.96 ;
		RECT	0 104.26 0.32 105.045 ;
		RECT	0 106.335 0.32 106.84 ;
		RECT	0 107.14 0.32 107.925 ;
		RECT	0 109.215 0.32 109.72 ;
		RECT	0 110.02 0.32 110.805 ;
		RECT	0 112.095 0.32 112.6 ;
		RECT	0 112.9 0.32 113.685 ;
		RECT	0 114.975 0.32 115.48 ;
		RECT	0 115.78 0.32 116.565 ;
		RECT	0 117.855 0.32 118.36 ;
		RECT	0 118.66 0.32 119.445 ;
		RECT	0 120.735 0.32 121.24 ;
		RECT	0 121.54 0.32 122.325 ;
		RECT	0 123.615 0.32 124.12 ;
		RECT	0 124.42 0.32 125.205 ;
		RECT	0 126.495 0.32 127 ;
		RECT	0 127.3 0.32 128.085 ;
		RECT	0 129.375 0.32 129.88 ;
		RECT	0 130.18 0.32 130.965 ;
		RECT	0 132.255 0.32 132.76 ;
		RECT	0 133.06 0.32 133.845 ;
		RECT	0 135.135 0.32 135.64 ;
		RECT	0 135.94 0.32 136.725 ;
		RECT	0 138.015 0.32 138.52 ;
		RECT	0 138.82 0.32 139.605 ;
		RECT	0 140.895 0.32 141.4 ;
		RECT	0 141.7 0.32 142.485 ;
		RECT	0 143.775 0.32 144.28 ;
		RECT	0 144.58 0.32 145.365 ;
		RECT	0 146.655 0.32 147.16 ;
		RECT	0 147.46 0.32 148.245 ;
		RECT	0 149.535 0.32 150.04 ;
		RECT	0 150.34 0.32 151.125 ;
		RECT	0 152.415 0.32 152.92 ;
		RECT	0 153.22 0.32 154.005 ;
		RECT	0 155.295 0.32 155.8 ;
		RECT	0 156.1 0.32 156.885 ;
		RECT	0 158.175 0.32 158.68 ;
		RECT	0 158.98 0.32 159.765 ;
		RECT	0 161.055 0.32 161.56 ;
		RECT	0 161.86 0.32 162.645 ;
		RECT	0 163.935 0.32 164.44 ;
		RECT	0 164.74 0.32 165.525 ;
		RECT	0 166.815 0.32 167.32 ;
		RECT	0 167.62 0.32 168.405 ;
		RECT	0 169.695 0.32 170.2 ;
		RECT	0 170.5 0.32 171.285 ;
		RECT	0 172.575 0.32 173.08 ;
		RECT	0 173.38 0.32 174.165 ;
		RECT	0 175.455 0.32 175.96 ;
		RECT	0 176.26 0.32 177.045 ;
		RECT	0 178.335 0.32 178.84 ;
		RECT	0 179.14 0.32 179.925 ;
		RECT	0 181.215 0.32 181.72 ;
		RECT	0 182.02 0.32 182.805 ;
		RECT	0 184.095 0.32 184.6 ;
		RECT	0 184.9 0.32 187 ;
		RECT	0 187.3 0.32 187.35 ;
		RECT	0 187.65 0.32 188.01 ;
		RECT	0 188.71 0.32 190.35 ;
		RECT	0 190.955 0.32 191.17 ;
		RECT	0 191.47 0.32 191.575 ;
		RECT	0 191.875 0.32 193.685 ;
		RECT	0 193.985 0.32 194.2 ;
		RECT	0 194.5 0.32 194.605 ;
		RECT	0 194.905 0.32 196.745 ;
		RECT	0 197.045 0.32 197.23 ;
		RECT	0 197.53 0.32 197.635 ;
		RECT	0 197.935 0.32 198.03 ;
		RECT	0 198.33 0.32 198.4 ;
		RECT	0 198.7 0.32 198.775 ;
		RECT	0 199.075 0.32 199.26 ;
		RECT	0 199.97 0.32 201.405 ;
		RECT	0 202.105 0.32 202.29 ;
		RECT	0 202.875 0.32 205.8 ;
		RECT	0 206.5 0.32 206.97 ;
		RECT	0 207.27 0.32 208.635 ;
		RECT	0 208.935 0.32 212.725 ;
		RECT	0 213.26 0.32 213.45 ;
		RECT	0 213.75 0.32 213.825 ;
		RECT	0 214.125 0.32 214.205 ;
		RECT	0 214.505 0.32 215.205 ;
		RECT	0 215.505 0.32 215.995 ;
		RECT	0 216.295 0.32 216.48 ;
		RECT	0 216.78 0.32 216.885 ;
		RECT	0 217.185 0.32 217.65 ;
		RECT	0 217.95 0.32 218.025 ;
		RECT	0 218.325 0.32 218.48 ;
		RECT	0 218.98 0.32 220.225 ;
		RECT	0 220.525 0.32 220.65 ;
		RECT	0 221.16 0.32 221.54 ;
		RECT	0 221.84 0.32 223.68 ;
		RECT	0 223.98 0.32 224.085 ;
		RECT	0 224.385 0.32 224.57 ;
		RECT	0 225.125 0.32 225.6 ;
		RECT	0 225.9 0.32 228.21 ;
		RECT	0 228.51 0.32 228.605 ;
		RECT	0 228.905 0.32 229.15 ;
		RECT	0 229.45 0.32 229.96 ;
		RECT	0 230.26 0.32 230.765 ;
		RECT	0 232.055 0.32 232.84 ;
		RECT	0 233.14 0.32 233.645 ;
		RECT	0 234.935 0.32 235.72 ;
		RECT	0 236.02 0.32 236.525 ;
		RECT	0 237.815 0.32 238.6 ;
		RECT	0 238.9 0.32 239.405 ;
		RECT	0 240.695 0.32 241.48 ;
		RECT	0 241.78 0.32 242.285 ;
		RECT	0 243.575 0.32 244.36 ;
		RECT	0 244.66 0.32 245.165 ;
		RECT	0 246.455 0.32 247.24 ;
		RECT	0 247.54 0.32 248.045 ;
		RECT	0 249.335 0.32 250.12 ;
		RECT	0 250.42 0.32 250.925 ;
		RECT	0 252.215 0.32 253 ;
		RECT	0 253.3 0.32 253.805 ;
		RECT	0 255.095 0.32 255.88 ;
		RECT	0 256.18 0.32 256.685 ;
		RECT	0 257.975 0.32 258.76 ;
		RECT	0 259.06 0.32 259.565 ;
		RECT	0 260.855 0.32 261.64 ;
		RECT	0 261.94 0.32 262.445 ;
		RECT	0 263.735 0.32 264.52 ;
		RECT	0 264.82 0.32 265.325 ;
		RECT	0 266.615 0.32 267.4 ;
		RECT	0 267.7 0.32 268.205 ;
		RECT	0 269.495 0.32 270.28 ;
		RECT	0 270.58 0.32 271.085 ;
		RECT	0 272.375 0.32 273.16 ;
		RECT	0 273.46 0.32 273.965 ;
		RECT	0 275.255 0.32 276.04 ;
		RECT	0 276.34 0.32 276.845 ;
		RECT	0 278.135 0.32 278.92 ;
		RECT	0 279.22 0.32 279.725 ;
		RECT	0 281.015 0.32 281.8 ;
		RECT	0 282.1 0.32 282.605 ;
		RECT	0 283.895 0.32 284.68 ;
		RECT	0 284.98 0.32 285.485 ;
		RECT	0 286.775 0.32 287.56 ;
		RECT	0 287.86 0.32 288.365 ;
		RECT	0 289.655 0.32 290.44 ;
		RECT	0 290.74 0.32 291.245 ;
		RECT	0 292.535 0.32 293.32 ;
		RECT	0 293.62 0.32 294.125 ;
		RECT	0 295.415 0.32 296.2 ;
		RECT	0 296.5 0.32 297.005 ;
		RECT	0 298.295 0.32 299.08 ;
		RECT	0 299.38 0.32 299.885 ;
		RECT	0 301.175 0.32 301.96 ;
		RECT	0 302.26 0.32 302.765 ;
		RECT	0 304.055 0.32 304.84 ;
		RECT	0 305.14 0.32 305.645 ;
		RECT	0 306.935 0.32 307.72 ;
		RECT	0 308.02 0.32 308.525 ;
		RECT	0 309.815 0.32 310.6 ;
		RECT	0 310.9 0.32 311.405 ;
		RECT	0 312.695 0.32 313.48 ;
		RECT	0 313.78 0.32 314.285 ;
		RECT	0 315.575 0.32 316.36 ;
		RECT	0 316.66 0.32 317.165 ;
		RECT	0 318.455 0.32 319.24 ;
		RECT	0 319.54 0.32 320.045 ;
		RECT	0 321.335 0.32 322.12 ;
		RECT	0 322.42 0.32 322.925 ;
		RECT	0 324.215 0.32 325 ;
		RECT	0 325.3 0.32 325.805 ;
		RECT	0 327.095 0.32 327.88 ;
		RECT	0 328.18 0.32 328.685 ;
		RECT	0 329.975 0.32 330.76 ;
		RECT	0 331.06 0.32 331.565 ;
		RECT	0 332.855 0.32 333.64 ;
		RECT	0 333.94 0.32 334.445 ;
		RECT	0 335.735 0.32 336.52 ;
		RECT	0 336.82 0.32 337.325 ;
		RECT	0 338.615 0.32 339.4 ;
		RECT	0 339.7 0.32 340.205 ;
		RECT	0 341.495 0.32 342.28 ;
		RECT	0 342.58 0.32 343.085 ;
		RECT	0 344.375 0.32 345.16 ;
		RECT	0 345.46 0.32 345.965 ;
		RECT	0 347.255 0.32 348.04 ;
		RECT	0 348.34 0.32 348.845 ;
		RECT	0 350.135 0.32 350.92 ;
		RECT	0 351.22 0.32 351.725 ;
		RECT	0 353.015 0.32 353.8 ;
		RECT	0 354.1 0.32 354.605 ;
		RECT	0 355.895 0.32 356.68 ;
		RECT	0 356.98 0.32 357.485 ;
		RECT	0 358.775 0.32 359.56 ;
		RECT	0 359.86 0.32 360.365 ;
		RECT	0 361.655 0.32 362.44 ;
		RECT	0 362.74 0.32 363.245 ;
		RECT	0 364.535 0.32 365.32 ;
		RECT	0 365.62 0.32 366.125 ;
		RECT	0 367.415 0.32 368.2 ;
		RECT	0 368.5 0.32 369.005 ;
		RECT	0 370.295 0.32 371.08 ;
		RECT	0 371.38 0.32 371.885 ;
		RECT	0 373.175 0.32 373.96 ;
		RECT	0 374.26 0.32 374.765 ;
		RECT	0 376.055 0.32 376.84 ;
		RECT	0 377.14 0.32 377.645 ;
		RECT	0 378.935 0.32 379.72 ;
		RECT	0 380.02 0.32 380.525 ;
		RECT	0 381.815 0.32 382.6 ;
		RECT	0 382.9 0.32 383.405 ;
		RECT	0 384.695 0.32 385.48 ;
		RECT	0 385.78 0.32 386.285 ;
		RECT	0 387.575 0.32 388.36 ;
		RECT	0 388.66 0.32 389.165 ;
		RECT	0 390.455 0.32 391.24 ;
		RECT	0 391.54 0.32 392.045 ;
		RECT	0 393.335 0.32 394.12 ;
		RECT	0 394.42 0.32 394.925 ;
		RECT	0 396.215 0.32 397 ;
		RECT	0 397.3 0.32 397.805 ;
		RECT	0 399.095 0.32 399.88 ;
		RECT	0 400.18 0.32 400.685 ;
		RECT	0 401.975 0.32 402.76 ;
		RECT	0 403.06 0.32 403.565 ;
		RECT	0 404.855 0.32 405.64 ;
		RECT	0 405.94 0.32 406.445 ;
		RECT	0 407.735 0.32 408.52 ;
		RECT	0 408.82 0.32 409.325 ;
		RECT	0 410.615 0.32 411.4 ;
		RECT	0 411.7 0.32 412.205 ;
		RECT	0 413.495 0.32 414.3 ;
		RECT	20.845 0 21.165 414.86 ;
		RECT	0.32 0 20.845 0.35 ;
		RECT	0.32 414.51 20.845 414.86 ;
		LAYER	M3 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 20.845 414.51 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 2.655 0.32 3.16 ;
		RECT	0 3.46 0.32 4.245 ;
		RECT	0 5.535 0.32 6.04 ;
		RECT	0 6.34 0.32 7.125 ;
		RECT	0 8.415 0.32 8.92 ;
		RECT	0 9.22 0.32 10.005 ;
		RECT	0 11.295 0.32 11.8 ;
		RECT	0 12.1 0.32 12.885 ;
		RECT	0 14.175 0.32 14.68 ;
		RECT	0 14.98 0.32 15.765 ;
		RECT	0 17.055 0.32 17.56 ;
		RECT	0 17.86 0.32 18.645 ;
		RECT	0 19.935 0.32 20.44 ;
		RECT	0 20.74 0.32 21.525 ;
		RECT	0 22.815 0.32 23.32 ;
		RECT	0 23.62 0.32 24.405 ;
		RECT	0 25.695 0.32 26.2 ;
		RECT	0 26.5 0.32 27.285 ;
		RECT	0 28.575 0.32 29.08 ;
		RECT	0 29.38 0.32 30.165 ;
		RECT	0 31.455 0.32 31.96 ;
		RECT	0 32.26 0.32 33.045 ;
		RECT	0 34.335 0.32 34.84 ;
		RECT	0 35.14 0.32 35.925 ;
		RECT	0 37.215 0.32 37.72 ;
		RECT	0 38.02 0.32 38.805 ;
		RECT	0 40.095 0.32 40.6 ;
		RECT	0 40.9 0.32 41.685 ;
		RECT	0 42.975 0.32 43.48 ;
		RECT	0 43.78 0.32 44.565 ;
		RECT	0 45.855 0.32 46.36 ;
		RECT	0 46.66 0.32 47.445 ;
		RECT	0 48.735 0.32 49.24 ;
		RECT	0 49.54 0.32 50.325 ;
		RECT	0 51.615 0.32 52.12 ;
		RECT	0 52.42 0.32 53.205 ;
		RECT	0 54.495 0.32 55 ;
		RECT	0 55.3 0.32 56.085 ;
		RECT	0 57.375 0.32 57.88 ;
		RECT	0 58.18 0.32 58.965 ;
		RECT	0 60.255 0.32 60.76 ;
		RECT	0 61.06 0.32 61.845 ;
		RECT	0 63.135 0.32 63.64 ;
		RECT	0 63.94 0.32 64.725 ;
		RECT	0 66.015 0.32 66.52 ;
		RECT	0 66.82 0.32 67.605 ;
		RECT	0 68.895 0.32 69.4 ;
		RECT	0 69.7 0.32 70.485 ;
		RECT	0 71.775 0.32 72.28 ;
		RECT	0 72.58 0.32 73.365 ;
		RECT	0 74.655 0.32 75.16 ;
		RECT	0 75.46 0.32 76.245 ;
		RECT	0 77.535 0.32 78.04 ;
		RECT	0 78.34 0.32 79.125 ;
		RECT	0 80.415 0.32 80.92 ;
		RECT	0 81.22 0.32 82.005 ;
		RECT	0 83.295 0.32 83.8 ;
		RECT	0 84.1 0.32 84.885 ;
		RECT	0 86.175 0.32 86.68 ;
		RECT	0 86.98 0.32 87.765 ;
		RECT	0 89.055 0.32 89.56 ;
		RECT	0 89.86 0.32 90.645 ;
		RECT	0 91.935 0.32 92.44 ;
		RECT	0 92.74 0.32 93.525 ;
		RECT	0 94.815 0.32 95.32 ;
		RECT	0 95.62 0.32 96.405 ;
		RECT	0 97.695 0.32 98.2 ;
		RECT	0 98.5 0.32 99.285 ;
		RECT	0 100.575 0.32 101.08 ;
		RECT	0 101.38 0.32 102.165 ;
		RECT	0 103.455 0.32 103.96 ;
		RECT	0 104.26 0.32 105.045 ;
		RECT	0 106.335 0.32 106.84 ;
		RECT	0 107.14 0.32 107.925 ;
		RECT	0 109.215 0.32 109.72 ;
		RECT	0 110.02 0.32 110.805 ;
		RECT	0 112.095 0.32 112.6 ;
		RECT	0 112.9 0.32 113.685 ;
		RECT	0 114.975 0.32 115.48 ;
		RECT	0 115.78 0.32 116.565 ;
		RECT	0 117.855 0.32 118.36 ;
		RECT	0 118.66 0.32 119.445 ;
		RECT	0 120.735 0.32 121.24 ;
		RECT	0 121.54 0.32 122.325 ;
		RECT	0 123.615 0.32 124.12 ;
		RECT	0 124.42 0.32 125.205 ;
		RECT	0 126.495 0.32 127 ;
		RECT	0 127.3 0.32 128.085 ;
		RECT	0 129.375 0.32 129.88 ;
		RECT	0 130.18 0.32 130.965 ;
		RECT	0 132.255 0.32 132.76 ;
		RECT	0 133.06 0.32 133.845 ;
		RECT	0 135.135 0.32 135.64 ;
		RECT	0 135.94 0.32 136.725 ;
		RECT	0 138.015 0.32 138.52 ;
		RECT	0 138.82 0.32 139.605 ;
		RECT	0 140.895 0.32 141.4 ;
		RECT	0 141.7 0.32 142.485 ;
		RECT	0 143.775 0.32 144.28 ;
		RECT	0 144.58 0.32 145.365 ;
		RECT	0 146.655 0.32 147.16 ;
		RECT	0 147.46 0.32 148.245 ;
		RECT	0 149.535 0.32 150.04 ;
		RECT	0 150.34 0.32 151.125 ;
		RECT	0 152.415 0.32 152.92 ;
		RECT	0 153.22 0.32 154.005 ;
		RECT	0 155.295 0.32 155.8 ;
		RECT	0 156.1 0.32 156.885 ;
		RECT	0 158.175 0.32 158.68 ;
		RECT	0 158.98 0.32 159.765 ;
		RECT	0 161.055 0.32 161.56 ;
		RECT	0 161.86 0.32 162.645 ;
		RECT	0 163.935 0.32 164.44 ;
		RECT	0 164.74 0.32 165.525 ;
		RECT	0 166.815 0.32 167.32 ;
		RECT	0 167.62 0.32 168.405 ;
		RECT	0 169.695 0.32 170.2 ;
		RECT	0 170.5 0.32 171.285 ;
		RECT	0 172.575 0.32 173.08 ;
		RECT	0 173.38 0.32 174.165 ;
		RECT	0 175.455 0.32 175.96 ;
		RECT	0 176.26 0.32 177.045 ;
		RECT	0 178.335 0.32 178.84 ;
		RECT	0 179.14 0.32 179.925 ;
		RECT	0 181.215 0.32 181.72 ;
		RECT	0 182.02 0.32 182.805 ;
		RECT	0 184.095 0.32 184.6 ;
		RECT	0 184.9 0.32 187 ;
		RECT	0 187.3 0.32 187.35 ;
		RECT	0 187.65 0.32 188.01 ;
		RECT	0 188.71 0.32 190.35 ;
		RECT	0 190.955 0.32 191.17 ;
		RECT	0 191.47 0.32 191.575 ;
		RECT	0 191.875 0.32 193.685 ;
		RECT	0 193.985 0.32 194.2 ;
		RECT	0 194.5 0.32 194.605 ;
		RECT	0 194.905 0.32 196.745 ;
		RECT	0 197.045 0.32 197.23 ;
		RECT	0 197.53 0.32 197.635 ;
		RECT	0 197.935 0.32 198.03 ;
		RECT	0 198.33 0.32 198.4 ;
		RECT	0 198.7 0.32 198.775 ;
		RECT	0 199.075 0.32 199.26 ;
		RECT	0 199.97 0.32 201.405 ;
		RECT	0 202.105 0.32 202.29 ;
		RECT	0 202.875 0.32 205.8 ;
		RECT	0 206.5 0.32 206.97 ;
		RECT	0 207.27 0.32 208.635 ;
		RECT	0 208.935 0.32 212.725 ;
		RECT	0 213.26 0.32 213.45 ;
		RECT	0 213.75 0.32 213.825 ;
		RECT	0 214.125 0.32 214.205 ;
		RECT	0 214.505 0.32 215.205 ;
		RECT	0 215.505 0.32 215.995 ;
		RECT	0 216.295 0.32 216.48 ;
		RECT	0 216.78 0.32 216.885 ;
		RECT	0 217.185 0.32 217.65 ;
		RECT	0 217.95 0.32 218.025 ;
		RECT	0 218.325 0.32 218.48 ;
		RECT	0 218.98 0.32 220.225 ;
		RECT	0 220.525 0.32 220.65 ;
		RECT	0 221.16 0.32 221.54 ;
		RECT	0 221.84 0.32 223.68 ;
		RECT	0 223.98 0.32 224.085 ;
		RECT	0 224.385 0.32 224.57 ;
		RECT	0 225.125 0.32 225.6 ;
		RECT	0 225.9 0.32 228.21 ;
		RECT	0 228.51 0.32 228.605 ;
		RECT	0 228.905 0.32 229.15 ;
		RECT	0 229.45 0.32 229.96 ;
		RECT	0 230.26 0.32 230.765 ;
		RECT	0 232.055 0.32 232.84 ;
		RECT	0 233.14 0.32 233.645 ;
		RECT	0 234.935 0.32 235.72 ;
		RECT	0 236.02 0.32 236.525 ;
		RECT	0 237.815 0.32 238.6 ;
		RECT	0 238.9 0.32 239.405 ;
		RECT	0 240.695 0.32 241.48 ;
		RECT	0 241.78 0.32 242.285 ;
		RECT	0 243.575 0.32 244.36 ;
		RECT	0 244.66 0.32 245.165 ;
		RECT	0 246.455 0.32 247.24 ;
		RECT	0 247.54 0.32 248.045 ;
		RECT	0 249.335 0.32 250.12 ;
		RECT	0 250.42 0.32 250.925 ;
		RECT	0 252.215 0.32 253 ;
		RECT	0 253.3 0.32 253.805 ;
		RECT	0 255.095 0.32 255.88 ;
		RECT	0 256.18 0.32 256.685 ;
		RECT	0 257.975 0.32 258.76 ;
		RECT	0 259.06 0.32 259.565 ;
		RECT	0 260.855 0.32 261.64 ;
		RECT	0 261.94 0.32 262.445 ;
		RECT	0 263.735 0.32 264.52 ;
		RECT	0 264.82 0.32 265.325 ;
		RECT	0 266.615 0.32 267.4 ;
		RECT	0 267.7 0.32 268.205 ;
		RECT	0 269.495 0.32 270.28 ;
		RECT	0 270.58 0.32 271.085 ;
		RECT	0 272.375 0.32 273.16 ;
		RECT	0 273.46 0.32 273.965 ;
		RECT	0 275.255 0.32 276.04 ;
		RECT	0 276.34 0.32 276.845 ;
		RECT	0 278.135 0.32 278.92 ;
		RECT	0 279.22 0.32 279.725 ;
		RECT	0 281.015 0.32 281.8 ;
		RECT	0 282.1 0.32 282.605 ;
		RECT	0 283.895 0.32 284.68 ;
		RECT	0 284.98 0.32 285.485 ;
		RECT	0 286.775 0.32 287.56 ;
		RECT	0 287.86 0.32 288.365 ;
		RECT	0 289.655 0.32 290.44 ;
		RECT	0 290.74 0.32 291.245 ;
		RECT	0 292.535 0.32 293.32 ;
		RECT	0 293.62 0.32 294.125 ;
		RECT	0 295.415 0.32 296.2 ;
		RECT	0 296.5 0.32 297.005 ;
		RECT	0 298.295 0.32 299.08 ;
		RECT	0 299.38 0.32 299.885 ;
		RECT	0 301.175 0.32 301.96 ;
		RECT	0 302.26 0.32 302.765 ;
		RECT	0 304.055 0.32 304.84 ;
		RECT	0 305.14 0.32 305.645 ;
		RECT	0 306.935 0.32 307.72 ;
		RECT	0 308.02 0.32 308.525 ;
		RECT	0 309.815 0.32 310.6 ;
		RECT	0 310.9 0.32 311.405 ;
		RECT	0 312.695 0.32 313.48 ;
		RECT	0 313.78 0.32 314.285 ;
		RECT	0 315.575 0.32 316.36 ;
		RECT	0 316.66 0.32 317.165 ;
		RECT	0 318.455 0.32 319.24 ;
		RECT	0 319.54 0.32 320.045 ;
		RECT	0 321.335 0.32 322.12 ;
		RECT	0 322.42 0.32 322.925 ;
		RECT	0 324.215 0.32 325 ;
		RECT	0 325.3 0.32 325.805 ;
		RECT	0 327.095 0.32 327.88 ;
		RECT	0 328.18 0.32 328.685 ;
		RECT	0 329.975 0.32 330.76 ;
		RECT	0 331.06 0.32 331.565 ;
		RECT	0 332.855 0.32 333.64 ;
		RECT	0 333.94 0.32 334.445 ;
		RECT	0 335.735 0.32 336.52 ;
		RECT	0 336.82 0.32 337.325 ;
		RECT	0 338.615 0.32 339.4 ;
		RECT	0 339.7 0.32 340.205 ;
		RECT	0 341.495 0.32 342.28 ;
		RECT	0 342.58 0.32 343.085 ;
		RECT	0 344.375 0.32 345.16 ;
		RECT	0 345.46 0.32 345.965 ;
		RECT	0 347.255 0.32 348.04 ;
		RECT	0 348.34 0.32 348.845 ;
		RECT	0 350.135 0.32 350.92 ;
		RECT	0 351.22 0.32 351.725 ;
		RECT	0 353.015 0.32 353.8 ;
		RECT	0 354.1 0.32 354.605 ;
		RECT	0 355.895 0.32 356.68 ;
		RECT	0 356.98 0.32 357.485 ;
		RECT	0 358.775 0.32 359.56 ;
		RECT	0 359.86 0.32 360.365 ;
		RECT	0 361.655 0.32 362.44 ;
		RECT	0 362.74 0.32 363.245 ;
		RECT	0 364.535 0.32 365.32 ;
		RECT	0 365.62 0.32 366.125 ;
		RECT	0 367.415 0.32 368.2 ;
		RECT	0 368.5 0.32 369.005 ;
		RECT	0 370.295 0.32 371.08 ;
		RECT	0 371.38 0.32 371.885 ;
		RECT	0 373.175 0.32 373.96 ;
		RECT	0 374.26 0.32 374.765 ;
		RECT	0 376.055 0.32 376.84 ;
		RECT	0 377.14 0.32 377.645 ;
		RECT	0 378.935 0.32 379.72 ;
		RECT	0 380.02 0.32 380.525 ;
		RECT	0 381.815 0.32 382.6 ;
		RECT	0 382.9 0.32 383.405 ;
		RECT	0 384.695 0.32 385.48 ;
		RECT	0 385.78 0.32 386.285 ;
		RECT	0 387.575 0.32 388.36 ;
		RECT	0 388.66 0.32 389.165 ;
		RECT	0 390.455 0.32 391.24 ;
		RECT	0 391.54 0.32 392.045 ;
		RECT	0 393.335 0.32 394.12 ;
		RECT	0 394.42 0.32 394.925 ;
		RECT	0 396.215 0.32 397 ;
		RECT	0 397.3 0.32 397.805 ;
		RECT	0 399.095 0.32 399.88 ;
		RECT	0 400.18 0.32 400.685 ;
		RECT	0 401.975 0.32 402.76 ;
		RECT	0 403.06 0.32 403.565 ;
		RECT	0 404.855 0.32 405.64 ;
		RECT	0 405.94 0.32 406.445 ;
		RECT	0 407.735 0.32 408.52 ;
		RECT	0 408.82 0.32 409.325 ;
		RECT	0 410.615 0.32 411.4 ;
		RECT	0 411.7 0.32 412.205 ;
		RECT	0 413.495 0.32 414.3 ;
		RECT	20.845 0 21.165 414.86 ;
		RECT	0.32 0 20.845 0.35 ;
		RECT	0.32 414.51 20.845 414.86 ;
		LAYER	M4 DESIGNRULEWIDTH 0.165 ;
		RECT	0.57 185.175 14.49 186.345 ;
		RECT	14.185 186.345 14.49 186.575 ;
		RECT	0.57 186.405 14.125 186.555 ;
		RECT	0.57 187.305 14.49 187.415 ;
		RECT	0.57 187.55 14.49 187.74 ;
		RECT	0.57 188.225 14.49 188.325 ;
		RECT	0.57 188.715 11.56 188.815 ;
		RECT	0.57 189.205 14.49 189.305 ;
		RECT	11.255 189.305 14.49 189.31 ;
		RECT	11.255 189.31 12.345 189.655 ;
		RECT	0.57 189.405 11.155 189.615 ;
		RECT	12.445 189.41 14.49 189.6 ;
		RECT	11.255 189.655 11.56 189.715 ;
		RECT	0.57 189.715 11.56 189.785 ;
		RECT	0.57 189.885 14.49 190.075 ;
		RECT	0.57 190.175 14.49 190.33 ;
		RECT	0.57 190.72 14.49 190.785 ;
		RECT	0.57 191.175 14.49 191.28 ;
		RECT	0.57 191.67 14.49 191.77 ;
		RECT	0.57 192.16 14.15 192.26 ;
		RECT	0.57 192.65 14.49 192.755 ;
		RECT	0.57 193.145 14.49 193.245 ;
		RECT	0.57 193.635 14.49 193.74 ;
		RECT	0.57 193.84 14.49 194.03 ;
		RECT	0.57 194.13 14.49 194.23 ;
		RECT	0.57 194.62 14.49 194.725 ;
		RECT	0.57 195.115 14.49 195.215 ;
		RECT	0.57 195.605 14.49 195.705 ;
		RECT	0.57 196.095 14.49 196.2 ;
		RECT	0.57 196.59 14.49 196.69 ;
		RECT	0.57 197.08 14.49 197.18 ;
		RECT	0.57 197.57 14.49 197.675 ;
		RECT	0.57 197.775 14.49 197.965 ;
		RECT	0.57 198.065 14.49 198.165 ;
		RECT	0.57 198.555 14.49 198.66 ;
		RECT	0.57 199.05 14.49 199.15 ;
		RECT	8.61 199.54 14.49 199.63 ;
		RECT	0.57 199.555 8.56 199.625 ;
		RECT	0.57 200.04 14.49 200.135 ;
		RECT	0.57 200.525 14.49 200.625 ;
		RECT	0.57 201.015 14.49 201.12 ;
		RECT	9.515 201.51 14.49 201.6 ;
		RECT	9.295 201.515 9.465 201.525 ;
		RECT	0.57 201.525 9.465 201.595 ;
		RECT	9.295 201.595 9.465 201.605 ;
		RECT	0.57 201.7 14.49 201.91 ;
		RECT	0.57 202.01 14.49 202.105 ;
		RECT	0.57 202.495 14.49 202.6 ;
		RECT	0.57 202.99 14.49 203.085 ;
		RECT	0.57 203.475 14.49 203.58 ;
		RECT	0.57 203.97 14.49 204.055 ;
		RECT	0.57 204.445 14.49 204.68 ;
		RECT	0.57 204.68 13.465 204.795 ;
		RECT	13.565 204.78 14.49 204.97 ;
		RECT	11.215 204.795 13.465 205.055 ;
		RECT	0.57 204.855 11.155 205.005 ;
		RECT	0.57 205.445 13.8 205.545 ;
		RECT	0.57 205.645 14.49 205.835 ;
		RECT	0.57 205.935 13.8 206.04 ;
		RECT	0.57 206.43 14.49 206.53 ;
		RECT	0.57 206.92 14.49 207.02 ;
		RECT	0.57 207.41 7.02 207.515 ;
		RECT	13.595 207.41 14.49 207.515 ;
		RECT	0.57 207.905 14.49 208.005 ;
		RECT	0.57 208.395 14.49 208.5 ;
		RECT	0.57 208.89 13.8 208.99 ;
		RECT	0.57 209.09 14.49 209.28 ;
		RECT	0.57 209.38 13.8 209.48 ;
		RECT	11.215 209.87 13.5 210.13 ;
		RECT	13.6 209.895 14.49 210.085 ;
		RECT	0.57 209.92 11.155 210.07 ;
		RECT	0.57 210.13 13.5 210.185 ;
		RECT	0.57 210.185 14.49 210.48 ;
		RECT	0.57 210.87 14.49 210.955 ;
		RECT	0.57 211.345 14.49 211.45 ;
		RECT	0.57 211.84 14.49 211.945 ;
		RECT	0.57 212.335 14.49 212.425 ;
		RECT	7.785 212.835 14.49 212.915 ;
		RECT	0.57 212.84 7.735 212.91 ;
		RECT	0.57 213.015 14.49 213.225 ;
		RECT	0.57 213.325 14.49 213.42 ;
		RECT	0.57 213.81 14.49 213.91 ;
		RECT	0.57 214.3 14.49 214.405 ;
		RECT	0.57 214.795 14.49 214.885 ;
		RECT	8.06 215.295 14.49 215.385 ;
		RECT	0.57 215.3 8.01 215.37 ;
		RECT	0.57 215.775 14.49 215.88 ;
		RECT	0.57 216.27 14.49 216.37 ;
		RECT	0.57 216.76 14.49 216.865 ;
		RECT	0.57 216.965 14.49 217.155 ;
		RECT	0.57 217.255 14.49 217.355 ;
		RECT	0.57 217.745 14.49 217.845 ;
		RECT	0.57 218.235 14.49 218.34 ;
		RECT	0.57 218.73 14.49 218.83 ;
		RECT	0.57 219.22 14.49 219.325 ;
		RECT	0.57 219.715 14.49 219.815 ;
		RECT	0.57 220.205 14.49 220.305 ;
		RECT	0.57 220.695 14.15 220.79 ;
		RECT	0.57 220.89 14.49 221.1 ;
		RECT	2.785 221.2 14.49 221.29 ;
		RECT	0.57 221.68 14.49 221.775 ;
		RECT	0.57 222.19 14.49 222.26 ;
		RECT	0.57 222.68 14.49 222.75 ;
		RECT	0.57 223.165 14.49 223.225 ;
		RECT	0.57 223.615 14.49 223.75 ;
		RECT	0.57 224.14 14.49 224.21 ;
		RECT	0.57 224.6 14.49 224.75 ;
		RECT	0.57 224.85 14.49 225.04 ;
		RECT	0.57 225.14 12.555 225.215 ;
		RECT	11.255 225.215 12.555 225.225 ;
		RECT	11.255 225.225 12.27 225.615 ;
		RECT	0.57 225.315 11.155 225.525 ;
		RECT	12.37 225.325 14.49 225.515 ;
		RECT	11.255 225.615 14.49 225.625 ;
		RECT	0.57 225.625 14.49 225.72 ;
		RECT	0.57 226.11 12.555 226.21 ;
		RECT	0.57 226.6 14.49 226.705 ;
		RECT	0.57 227.105 14.49 227.315 ;
		RECT	0.57 227.445 14.49 227.555 ;
		RECT	14.21 228.285 14.49 228.515 ;
		RECT	0.57 228.305 14.15 228.455 ;
		RECT	0.57 228.515 14.49 229.685 ;
		RECT	0.21 186.405 0.57 186.555 ;
		RECT	0.215 187.55 0.57 187.74 ;
		RECT	0.22 189.405 0.57 189.615 ;
		RECT	0.22 189.885 0.57 190.075 ;
		RECT	0.22 193.84 0.57 194.03 ;
		RECT	0.23 197.775 0.57 197.965 ;
		RECT	0.14 199.555 0.57 199.625 ;
		RECT	0.15 201.525 0.57 201.595 ;
		RECT	0.215 201.7 0.57 201.91 ;
		RECT	0.21 204.855 0.57 205.005 ;
		RECT	0.225 205.645 0.57 205.835 ;
		RECT	0.325 209.09 0.61 209.28 ;
		RECT	0.21 209.92 0.57 210.07 ;
		RECT	0.15 212.84 0.57 212.91 ;
		RECT	0.235 213.015 0.57 213.225 ;
		RECT	0.14 215.3 0.57 215.37 ;
		RECT	0.24 216.965 0.57 217.155 ;
		RECT	0.225 220.89 0.57 221.1 ;
		RECT	0.14 221.205 0.57 221.275 ;
		RECT	0.235 224.85 0.57 225.04 ;
		RECT	0.225 225.315 0.57 225.525 ;
		RECT	0.24 227.105 0.57 227.315 ;
		RECT	0.22 228.305 0.57 228.455 ;
		RECT	5.7 181.625 13.945 181.775 ;
		RECT	5.7 155.705 13.945 155.855 ;
		RECT	5.7 152.825 13.945 152.975 ;
		RECT	5.7 149.945 13.945 150.095 ;
		RECT	5.7 147.065 13.945 147.215 ;
		RECT	5.7 144.185 13.945 144.335 ;
		RECT	5.7 141.305 13.945 141.455 ;
		RECT	5.7 138.425 13.945 138.575 ;
		RECT	5.7 135.545 13.945 135.695 ;
		RECT	5.7 132.665 13.945 132.815 ;
		RECT	5.7 129.785 13.945 129.935 ;
		RECT	5.7 178.745 13.945 178.895 ;
		RECT	5.7 126.905 13.945 127.055 ;
		RECT	5.7 124.025 13.945 124.175 ;
		RECT	5.7 121.145 13.945 121.295 ;
		RECT	5.7 118.265 13.945 118.415 ;
		RECT	5.7 115.385 13.945 115.535 ;
		RECT	5.7 112.505 13.945 112.655 ;
		RECT	5.7 109.625 13.945 109.775 ;
		RECT	5.7 106.745 13.945 106.895 ;
		RECT	5.7 103.865 13.945 104.015 ;
		RECT	5.7 100.985 13.945 101.135 ;
		RECT	5.7 175.865 13.945 176.015 ;
		RECT	5.7 98.105 13.945 98.255 ;
		RECT	5.7 95.225 13.945 95.375 ;
		RECT	5.7 92.345 13.945 92.495 ;
		RECT	5.7 89.465 13.945 89.615 ;
		RECT	5.7 86.585 13.945 86.735 ;
		RECT	5.7 83.705 13.945 83.855 ;
		RECT	5.7 80.825 13.945 80.975 ;
		RECT	5.7 77.945 13.945 78.095 ;
		RECT	5.7 75.065 13.945 75.215 ;
		RECT	5.7 72.185 13.945 72.335 ;
		RECT	5.7 172.985 13.945 173.135 ;
		RECT	5.7 69.305 13.945 69.455 ;
		RECT	5.7 66.425 13.945 66.575 ;
		RECT	5.7 63.545 13.945 63.695 ;
		RECT	5.7 60.665 13.945 60.815 ;
		RECT	5.7 57.785 13.945 57.935 ;
		RECT	5.7 54.905 13.945 55.055 ;
		RECT	5.7 52.025 13.945 52.175 ;
		RECT	5.7 49.145 13.945 49.295 ;
		RECT	5.7 46.265 13.945 46.415 ;
		RECT	5.7 43.385 13.945 43.535 ;
		RECT	5.7 170.105 13.945 170.255 ;
		RECT	5.7 40.505 13.945 40.655 ;
		RECT	5.7 37.625 13.945 37.775 ;
		RECT	5.7 34.745 13.945 34.895 ;
		RECT	5.7 31.865 13.945 32.015 ;
		RECT	5.7 28.985 13.945 29.135 ;
		RECT	5.7 26.105 13.945 26.255 ;
		RECT	5.7 23.225 13.945 23.375 ;
		RECT	5.7 20.345 13.945 20.495 ;
		RECT	5.7 17.465 13.945 17.615 ;
		RECT	5.7 14.585 13.945 14.735 ;
		RECT	5.7 167.225 13.945 167.375 ;
		RECT	5.7 11.705 13.945 11.855 ;
		RECT	5.7 8.825 13.945 8.975 ;
		RECT	5.7 5.945 13.945 6.095 ;
		RECT	5.7 164.345 13.945 164.495 ;
		RECT	5.7 161.465 13.945 161.615 ;
		RECT	5.7 158.585 13.945 158.735 ;
		RECT	5.7 3.065 13.945 3.215 ;
		RECT	5.7 184.505 13.945 184.655 ;
		RECT	0.57 181.625 1.11 181.775 ;
		RECT	0.57 155.705 1.11 155.855 ;
		RECT	0.57 152.825 1.11 152.975 ;
		RECT	0.57 149.945 1.11 150.095 ;
		RECT	0.57 147.065 1.11 147.215 ;
		RECT	0.57 144.185 1.11 144.335 ;
		RECT	0.57 141.305 1.11 141.455 ;
		RECT	0.57 138.425 1.11 138.575 ;
		RECT	0.57 135.545 1.11 135.695 ;
		RECT	0.57 132.665 1.11 132.815 ;
		RECT	0.57 129.785 1.11 129.935 ;
		RECT	0.57 178.745 1.11 178.895 ;
		RECT	0.57 126.905 1.11 127.055 ;
		RECT	0.57 124.025 1.11 124.175 ;
		RECT	0.57 121.145 1.11 121.295 ;
		RECT	0.57 118.265 1.11 118.415 ;
		RECT	0.57 115.385 1.11 115.535 ;
		RECT	0.57 112.505 1.11 112.655 ;
		RECT	0.57 109.625 1.11 109.775 ;
		RECT	0.57 106.745 1.11 106.895 ;
		RECT	0.57 103.865 1.11 104.015 ;
		RECT	0.57 100.985 1.11 101.135 ;
		RECT	0.57 175.865 1.11 176.015 ;
		RECT	0.57 98.105 1.11 98.255 ;
		RECT	0.57 95.225 1.11 95.375 ;
		RECT	0.57 92.345 1.11 92.495 ;
		RECT	0.57 89.465 1.11 89.615 ;
		RECT	0.57 86.585 1.11 86.735 ;
		RECT	0.57 83.705 1.11 83.855 ;
		RECT	0.57 80.825 1.11 80.975 ;
		RECT	0.57 77.945 1.11 78.095 ;
		RECT	0.57 75.065 1.11 75.215 ;
		RECT	0.57 72.185 1.11 72.335 ;
		RECT	0.57 172.985 1.11 173.135 ;
		RECT	0.57 69.305 1.11 69.455 ;
		RECT	0.57 66.425 1.11 66.575 ;
		RECT	0.57 63.545 1.11 63.695 ;
		RECT	0.57 60.665 1.11 60.815 ;
		RECT	0.57 57.785 1.11 57.935 ;
		RECT	0.57 54.905 1.11 55.055 ;
		RECT	0.57 52.025 1.11 52.175 ;
		RECT	0.57 49.145 1.11 49.295 ;
		RECT	0.57 46.265 1.11 46.415 ;
		RECT	0.57 43.385 1.11 43.535 ;
		RECT	0.57 170.105 1.11 170.255 ;
		RECT	0.57 40.505 1.11 40.655 ;
		RECT	0.57 37.625 1.11 37.775 ;
		RECT	0.57 34.745 1.11 34.895 ;
		RECT	0.57 31.865 1.11 32.015 ;
		RECT	0.57 28.985 1.11 29.135 ;
		RECT	0.57 26.105 1.11 26.255 ;
		RECT	0.57 23.225 1.11 23.375 ;
		RECT	0.57 20.345 1.11 20.495 ;
		RECT	0.57 17.465 1.11 17.615 ;
		RECT	0.57 14.585 1.11 14.735 ;
		RECT	0.57 167.225 1.11 167.375 ;
		RECT	0.57 11.705 1.11 11.855 ;
		RECT	0.57 8.825 1.11 8.975 ;
		RECT	0.57 5.945 1.11 6.095 ;
		RECT	0.57 164.345 1.11 164.495 ;
		RECT	0.57 161.465 1.11 161.615 ;
		RECT	0.57 158.585 1.11 158.735 ;
		RECT	0.57 3.065 1.11 3.215 ;
		RECT	0.57 184.505 1.11 184.655 ;
		RECT	1.005 181.625 5.7 181.775 ;
		RECT	1.005 155.705 5.7 155.855 ;
		RECT	1.005 152.825 5.7 152.975 ;
		RECT	1.005 149.945 5.7 150.095 ;
		RECT	1.005 147.065 5.7 147.215 ;
		RECT	1.005 144.185 5.7 144.335 ;
		RECT	1.005 141.305 5.7 141.455 ;
		RECT	1.005 138.425 5.7 138.575 ;
		RECT	1.005 135.545 5.7 135.695 ;
		RECT	1.005 132.665 5.7 132.815 ;
		RECT	1.005 129.785 5.7 129.935 ;
		RECT	1.005 178.745 5.7 178.895 ;
		RECT	1.005 126.905 5.7 127.055 ;
		RECT	1.005 124.025 5.7 124.175 ;
		RECT	1.005 121.145 5.7 121.295 ;
		RECT	1.005 118.265 5.7 118.415 ;
		RECT	1.005 115.385 5.7 115.535 ;
		RECT	1.005 112.505 5.7 112.655 ;
		RECT	1.005 109.625 5.7 109.775 ;
		RECT	1.005 106.745 5.7 106.895 ;
		RECT	1.005 103.865 5.7 104.015 ;
		RECT	1.005 100.985 5.7 101.135 ;
		RECT	1.005 175.865 5.7 176.015 ;
		RECT	1.005 98.105 5.7 98.255 ;
		RECT	1.005 95.225 5.7 95.375 ;
		RECT	1.005 92.345 5.7 92.495 ;
		RECT	1.005 89.465 5.7 89.615 ;
		RECT	1.005 86.585 5.7 86.735 ;
		RECT	1.005 83.705 5.7 83.855 ;
		RECT	1.005 80.825 5.7 80.975 ;
		RECT	1.005 77.945 5.7 78.095 ;
		RECT	1.005 75.065 5.7 75.215 ;
		RECT	1.005 72.185 5.7 72.335 ;
		RECT	1.005 172.985 5.7 173.135 ;
		RECT	1.005 69.305 5.7 69.455 ;
		RECT	1.005 66.425 5.7 66.575 ;
		RECT	1.005 63.545 5.7 63.695 ;
		RECT	1.005 60.665 5.7 60.815 ;
		RECT	1.005 57.785 5.7 57.935 ;
		RECT	1.005 54.905 5.7 55.055 ;
		RECT	1.005 52.025 5.7 52.175 ;
		RECT	1.005 49.145 5.7 49.295 ;
		RECT	1.005 46.265 5.7 46.415 ;
		RECT	1.005 43.385 5.7 43.535 ;
		RECT	1.005 170.105 5.7 170.255 ;
		RECT	1.005 40.505 5.7 40.655 ;
		RECT	1.005 37.625 5.7 37.775 ;
		RECT	1.005 34.745 5.7 34.895 ;
		RECT	1.005 31.865 5.7 32.015 ;
		RECT	1.005 28.985 5.7 29.135 ;
		RECT	1.005 26.105 5.7 26.255 ;
		RECT	1.005 23.225 5.7 23.375 ;
		RECT	1.005 20.345 5.7 20.495 ;
		RECT	1.005 17.465 5.7 17.615 ;
		RECT	1.005 14.585 5.7 14.735 ;
		RECT	1.005 167.225 5.7 167.375 ;
		RECT	1.005 11.705 5.7 11.855 ;
		RECT	1.005 8.825 5.7 8.975 ;
		RECT	1.005 5.945 5.7 6.095 ;
		RECT	1.005 164.345 5.7 164.495 ;
		RECT	1.005 161.465 5.7 161.615 ;
		RECT	1.005 158.585 5.7 158.735 ;
		RECT	1.005 3.065 5.7 3.215 ;
		RECT	1.005 184.505 5.7 184.655 ;
		RECT	0.255 184.505 0.57 184.655 ;
		RECT	0.255 181.625 0.57 181.775 ;
		RECT	0.255 155.705 0.57 155.855 ;
		RECT	0.255 152.825 0.57 152.975 ;
		RECT	0.255 149.945 0.57 150.095 ;
		RECT	0.255 147.065 0.57 147.215 ;
		RECT	0.255 144.185 0.57 144.335 ;
		RECT	0.255 141.305 0.57 141.455 ;
		RECT	0.255 138.425 0.57 138.575 ;
		RECT	0.255 135.545 0.57 135.695 ;
		RECT	0.255 132.665 0.57 132.815 ;
		RECT	0.255 129.785 0.57 129.935 ;
		RECT	0.255 178.745 0.57 178.895 ;
		RECT	0.255 126.905 0.57 127.055 ;
		RECT	0.255 124.025 0.57 124.175 ;
		RECT	0.255 121.145 0.57 121.295 ;
		RECT	0.255 118.265 0.57 118.415 ;
		RECT	0.255 115.385 0.57 115.535 ;
		RECT	0.255 112.505 0.57 112.655 ;
		RECT	0.255 109.625 0.57 109.775 ;
		RECT	0.255 106.745 0.57 106.895 ;
		RECT	0.255 103.865 0.57 104.015 ;
		RECT	0.255 100.985 0.57 101.135 ;
		RECT	0.255 175.865 0.57 176.015 ;
		RECT	0.255 98.105 0.57 98.255 ;
		RECT	0.255 95.225 0.57 95.375 ;
		RECT	0.255 92.345 0.57 92.495 ;
		RECT	0.255 89.465 0.57 89.615 ;
		RECT	0.255 86.585 0.57 86.735 ;
		RECT	0.255 83.705 0.57 83.855 ;
		RECT	0.255 80.825 0.57 80.975 ;
		RECT	0.255 77.945 0.57 78.095 ;
		RECT	0.255 75.065 0.57 75.215 ;
		RECT	0.255 72.185 0.57 72.335 ;
		RECT	0.255 172.985 0.57 173.135 ;
		RECT	0.255 69.305 0.57 69.455 ;
		RECT	0.255 66.425 0.57 66.575 ;
		RECT	0.255 63.545 0.57 63.695 ;
		RECT	0.255 60.665 0.57 60.815 ;
		RECT	0.255 57.785 0.57 57.935 ;
		RECT	0.255 54.905 0.57 55.055 ;
		RECT	0.255 52.025 0.57 52.175 ;
		RECT	0.255 49.145 0.57 49.295 ;
		RECT	0.255 46.265 0.57 46.415 ;
		RECT	0.255 43.385 0.57 43.535 ;
		RECT	0.255 170.105 0.57 170.255 ;
		RECT	0.255 40.505 0.57 40.655 ;
		RECT	0.255 37.625 0.57 37.775 ;
		RECT	0.255 34.745 0.57 34.895 ;
		RECT	0.255 31.865 0.57 32.015 ;
		RECT	0.255 28.985 0.57 29.135 ;
		RECT	0.255 26.105 0.57 26.255 ;
		RECT	0.255 23.225 0.57 23.375 ;
		RECT	0.255 20.345 0.57 20.495 ;
		RECT	0.255 17.465 0.57 17.615 ;
		RECT	0.255 14.585 0.57 14.735 ;
		RECT	0.255 167.225 0.57 167.375 ;
		RECT	0.255 11.705 0.57 11.855 ;
		RECT	0.255 8.825 0.57 8.975 ;
		RECT	0.255 5.945 0.57 6.095 ;
		RECT	0.255 3.065 0.57 3.215 ;
		RECT	0.255 164.345 0.57 164.495 ;
		RECT	0.255 161.465 0.57 161.615 ;
		RECT	0.255 158.585 0.57 158.735 ;
		RECT	5.7 233.085 13.945 233.235 ;
		RECT	5.7 259.005 13.945 259.155 ;
		RECT	5.7 261.885 13.945 262.035 ;
		RECT	5.7 264.765 13.945 264.915 ;
		RECT	5.7 267.645 13.945 267.795 ;
		RECT	5.7 270.525 13.945 270.675 ;
		RECT	5.7 273.405 13.945 273.555 ;
		RECT	5.7 276.285 13.945 276.435 ;
		RECT	5.7 279.165 13.945 279.315 ;
		RECT	5.7 282.045 13.945 282.195 ;
		RECT	5.7 284.925 13.945 285.075 ;
		RECT	5.7 235.965 13.945 236.115 ;
		RECT	5.7 287.805 13.945 287.955 ;
		RECT	5.7 290.685 13.945 290.835 ;
		RECT	5.7 293.565 13.945 293.715 ;
		RECT	5.7 296.445 13.945 296.595 ;
		RECT	5.7 299.325 13.945 299.475 ;
		RECT	5.7 302.205 13.945 302.355 ;
		RECT	5.7 305.085 13.945 305.235 ;
		RECT	5.7 307.965 13.945 308.115 ;
		RECT	5.7 310.845 13.945 310.995 ;
		RECT	5.7 313.725 13.945 313.875 ;
		RECT	5.7 238.845 13.945 238.995 ;
		RECT	5.7 316.605 13.945 316.755 ;
		RECT	5.7 319.485 13.945 319.635 ;
		RECT	5.7 322.365 13.945 322.515 ;
		RECT	5.7 325.245 13.945 325.395 ;
		RECT	5.7 328.125 13.945 328.275 ;
		RECT	5.7 331.005 13.945 331.155 ;
		RECT	5.7 333.885 13.945 334.035 ;
		RECT	5.7 336.765 13.945 336.915 ;
		RECT	5.7 339.645 13.945 339.795 ;
		RECT	5.7 342.525 13.945 342.675 ;
		RECT	5.7 241.725 13.945 241.875 ;
		RECT	5.7 345.405 13.945 345.555 ;
		RECT	5.7 348.285 13.945 348.435 ;
		RECT	5.7 351.165 13.945 351.315 ;
		RECT	5.7 354.045 13.945 354.195 ;
		RECT	5.7 356.925 13.945 357.075 ;
		RECT	5.7 359.805 13.945 359.955 ;
		RECT	5.7 362.685 13.945 362.835 ;
		RECT	5.7 365.565 13.945 365.715 ;
		RECT	5.7 368.445 13.945 368.595 ;
		RECT	5.7 371.325 13.945 371.475 ;
		RECT	5.7 244.605 13.945 244.755 ;
		RECT	5.7 374.205 13.945 374.355 ;
		RECT	5.7 377.085 13.945 377.235 ;
		RECT	5.7 379.965 13.945 380.115 ;
		RECT	5.7 382.845 13.945 382.995 ;
		RECT	5.7 385.725 13.945 385.875 ;
		RECT	5.7 388.605 13.945 388.755 ;
		RECT	5.7 391.485 13.945 391.635 ;
		RECT	5.7 394.365 13.945 394.515 ;
		RECT	5.7 397.245 13.945 397.395 ;
		RECT	5.7 400.125 13.945 400.275 ;
		RECT	5.7 247.485 13.945 247.635 ;
		RECT	5.7 403.005 13.945 403.155 ;
		RECT	5.7 405.885 13.945 406.035 ;
		RECT	5.7 408.765 13.945 408.915 ;
		RECT	5.7 250.365 13.945 250.515 ;
		RECT	5.7 253.245 13.945 253.395 ;
		RECT	5.7 256.125 13.945 256.275 ;
		RECT	5.7 411.645 13.945 411.795 ;
		RECT	5.7 230.205 13.945 230.355 ;
		RECT	0.57 233.085 1.11 233.235 ;
		RECT	0.57 259.005 1.11 259.155 ;
		RECT	0.57 261.885 1.11 262.035 ;
		RECT	0.57 264.765 1.11 264.915 ;
		RECT	0.57 267.645 1.11 267.795 ;
		RECT	0.57 270.525 1.11 270.675 ;
		RECT	0.57 273.405 1.11 273.555 ;
		RECT	0.57 276.285 1.11 276.435 ;
		RECT	0.57 279.165 1.11 279.315 ;
		RECT	0.57 282.045 1.11 282.195 ;
		RECT	0.57 284.925 1.11 285.075 ;
		RECT	0.57 235.965 1.11 236.115 ;
		RECT	0.57 287.805 1.11 287.955 ;
		RECT	0.57 290.685 1.11 290.835 ;
		RECT	0.57 293.565 1.11 293.715 ;
		RECT	0.57 296.445 1.11 296.595 ;
		RECT	0.57 299.325 1.11 299.475 ;
		RECT	0.57 302.205 1.11 302.355 ;
		RECT	0.57 305.085 1.11 305.235 ;
		RECT	0.57 307.965 1.11 308.115 ;
		RECT	0.57 310.845 1.11 310.995 ;
		RECT	0.57 313.725 1.11 313.875 ;
		RECT	0.57 238.845 1.11 238.995 ;
		RECT	0.57 316.605 1.11 316.755 ;
		RECT	0.57 319.485 1.11 319.635 ;
		RECT	0.57 322.365 1.11 322.515 ;
		RECT	0.57 325.245 1.11 325.395 ;
		RECT	0.57 328.125 1.11 328.275 ;
		RECT	0.57 331.005 1.11 331.155 ;
		RECT	0.57 333.885 1.11 334.035 ;
		RECT	0.57 336.765 1.11 336.915 ;
		RECT	0.57 339.645 1.11 339.795 ;
		RECT	0.57 342.525 1.11 342.675 ;
		RECT	0.57 241.725 1.11 241.875 ;
		RECT	0.57 345.405 1.11 345.555 ;
		RECT	0.57 348.285 1.11 348.435 ;
		RECT	0.57 351.165 1.11 351.315 ;
		RECT	0.57 354.045 1.11 354.195 ;
		RECT	0.57 356.925 1.11 357.075 ;
		RECT	0.57 359.805 1.11 359.955 ;
		RECT	0.57 362.685 1.11 362.835 ;
		RECT	0.57 365.565 1.11 365.715 ;
		RECT	0.57 368.445 1.11 368.595 ;
		RECT	0.57 371.325 1.11 371.475 ;
		RECT	0.57 244.605 1.11 244.755 ;
		RECT	0.57 374.205 1.11 374.355 ;
		RECT	0.57 377.085 1.11 377.235 ;
		RECT	0.57 379.965 1.11 380.115 ;
		RECT	0.57 382.845 1.11 382.995 ;
		RECT	0.57 385.725 1.11 385.875 ;
		RECT	0.57 388.605 1.11 388.755 ;
		RECT	0.57 391.485 1.11 391.635 ;
		RECT	0.57 394.365 1.11 394.515 ;
		RECT	0.57 397.245 1.11 397.395 ;
		RECT	0.57 400.125 1.11 400.275 ;
		RECT	0.57 247.485 1.11 247.635 ;
		RECT	0.57 403.005 1.11 403.155 ;
		RECT	0.57 405.885 1.11 406.035 ;
		RECT	0.57 408.765 1.11 408.915 ;
		RECT	0.57 250.365 1.11 250.515 ;
		RECT	0.57 253.245 1.11 253.395 ;
		RECT	0.57 256.125 1.11 256.275 ;
		RECT	0.57 411.645 1.11 411.795 ;
		RECT	0.57 230.205 1.11 230.355 ;
		RECT	1.005 233.085 5.7 233.235 ;
		RECT	1.005 259.005 5.7 259.155 ;
		RECT	1.005 261.885 5.7 262.035 ;
		RECT	1.005 264.765 5.7 264.915 ;
		RECT	1.005 267.645 5.7 267.795 ;
		RECT	1.005 270.525 5.7 270.675 ;
		RECT	1.005 273.405 5.7 273.555 ;
		RECT	1.005 276.285 5.7 276.435 ;
		RECT	1.005 279.165 5.7 279.315 ;
		RECT	1.005 282.045 5.7 282.195 ;
		RECT	1.005 284.925 5.7 285.075 ;
		RECT	1.005 235.965 5.7 236.115 ;
		RECT	1.005 287.805 5.7 287.955 ;
		RECT	1.005 290.685 5.7 290.835 ;
		RECT	1.005 293.565 5.7 293.715 ;
		RECT	1.005 296.445 5.7 296.595 ;
		RECT	1.005 299.325 5.7 299.475 ;
		RECT	1.005 302.205 5.7 302.355 ;
		RECT	1.005 305.085 5.7 305.235 ;
		RECT	1.005 307.965 5.7 308.115 ;
		RECT	1.005 310.845 5.7 310.995 ;
		RECT	1.005 313.725 5.7 313.875 ;
		RECT	1.005 238.845 5.7 238.995 ;
		RECT	1.005 316.605 5.7 316.755 ;
		RECT	1.005 319.485 5.7 319.635 ;
		RECT	1.005 322.365 5.7 322.515 ;
		RECT	1.005 325.245 5.7 325.395 ;
		RECT	1.005 328.125 5.7 328.275 ;
		RECT	1.005 331.005 5.7 331.155 ;
		RECT	1.005 333.885 5.7 334.035 ;
		RECT	1.005 336.765 5.7 336.915 ;
		RECT	1.005 339.645 5.7 339.795 ;
		RECT	1.005 342.525 5.7 342.675 ;
		RECT	1.005 241.725 5.7 241.875 ;
		RECT	1.005 345.405 5.7 345.555 ;
		RECT	1.005 348.285 5.7 348.435 ;
		RECT	1.005 351.165 5.7 351.315 ;
		RECT	1.005 354.045 5.7 354.195 ;
		RECT	1.005 356.925 5.7 357.075 ;
		RECT	1.005 359.805 5.7 359.955 ;
		RECT	1.005 362.685 5.7 362.835 ;
		RECT	1.005 365.565 5.7 365.715 ;
		RECT	1.005 368.445 5.7 368.595 ;
		RECT	1.005 371.325 5.7 371.475 ;
		RECT	1.005 244.605 5.7 244.755 ;
		RECT	1.005 374.205 5.7 374.355 ;
		RECT	1.005 377.085 5.7 377.235 ;
		RECT	1.005 379.965 5.7 380.115 ;
		RECT	1.005 382.845 5.7 382.995 ;
		RECT	1.005 385.725 5.7 385.875 ;
		RECT	1.005 388.605 5.7 388.755 ;
		RECT	1.005 391.485 5.7 391.635 ;
		RECT	1.005 394.365 5.7 394.515 ;
		RECT	1.005 397.245 5.7 397.395 ;
		RECT	1.005 400.125 5.7 400.275 ;
		RECT	1.005 247.485 5.7 247.635 ;
		RECT	1.005 403.005 5.7 403.155 ;
		RECT	1.005 405.885 5.7 406.035 ;
		RECT	1.005 408.765 5.7 408.915 ;
		RECT	1.005 250.365 5.7 250.515 ;
		RECT	1.005 253.245 5.7 253.395 ;
		RECT	1.005 256.125 5.7 256.275 ;
		RECT	1.005 411.645 5.7 411.795 ;
		RECT	1.005 230.205 5.7 230.355 ;
		RECT	0.255 230.205 0.57 230.355 ;
		RECT	0.255 233.085 0.57 233.235 ;
		RECT	0.255 259.005 0.57 259.155 ;
		RECT	0.255 261.885 0.57 262.035 ;
		RECT	0.255 264.765 0.57 264.915 ;
		RECT	0.255 267.645 0.57 267.795 ;
		RECT	0.255 270.525 0.57 270.675 ;
		RECT	0.255 273.405 0.57 273.555 ;
		RECT	0.255 276.285 0.57 276.435 ;
		RECT	0.255 279.165 0.57 279.315 ;
		RECT	0.255 282.045 0.57 282.195 ;
		RECT	0.255 284.925 0.57 285.075 ;
		RECT	0.255 235.965 0.57 236.115 ;
		RECT	0.255 287.805 0.57 287.955 ;
		RECT	0.255 290.685 0.57 290.835 ;
		RECT	0.255 293.565 0.57 293.715 ;
		RECT	0.255 296.445 0.57 296.595 ;
		RECT	0.255 299.325 0.57 299.475 ;
		RECT	0.255 302.205 0.57 302.355 ;
		RECT	0.255 305.085 0.57 305.235 ;
		RECT	0.255 307.965 0.57 308.115 ;
		RECT	0.255 310.845 0.57 310.995 ;
		RECT	0.255 313.725 0.57 313.875 ;
		RECT	0.255 238.845 0.57 238.995 ;
		RECT	0.255 316.605 0.57 316.755 ;
		RECT	0.255 319.485 0.57 319.635 ;
		RECT	0.255 322.365 0.57 322.515 ;
		RECT	0.255 325.245 0.57 325.395 ;
		RECT	0.255 328.125 0.57 328.275 ;
		RECT	0.255 331.005 0.57 331.155 ;
		RECT	0.255 333.885 0.57 334.035 ;
		RECT	0.255 336.765 0.57 336.915 ;
		RECT	0.255 339.645 0.57 339.795 ;
		RECT	0.255 342.525 0.57 342.675 ;
		RECT	0.255 241.725 0.57 241.875 ;
		RECT	0.255 345.405 0.57 345.555 ;
		RECT	0.255 348.285 0.57 348.435 ;
		RECT	0.255 351.165 0.57 351.315 ;
		RECT	0.255 354.045 0.57 354.195 ;
		RECT	0.255 356.925 0.57 357.075 ;
		RECT	0.255 359.805 0.57 359.955 ;
		RECT	0.255 362.685 0.57 362.835 ;
		RECT	0.255 365.565 0.57 365.715 ;
		RECT	0.255 368.445 0.57 368.595 ;
		RECT	0.255 371.325 0.57 371.475 ;
		RECT	0.255 244.605 0.57 244.755 ;
		RECT	0.255 374.205 0.57 374.355 ;
		RECT	0.255 377.085 0.57 377.235 ;
		RECT	0.255 379.965 0.57 380.115 ;
		RECT	0.255 382.845 0.57 382.995 ;
		RECT	0.255 385.725 0.57 385.875 ;
		RECT	0.255 388.605 0.57 388.755 ;
		RECT	0.255 391.485 0.57 391.635 ;
		RECT	0.255 394.365 0.57 394.515 ;
		RECT	0.255 397.245 0.57 397.395 ;
		RECT	0.255 400.125 0.57 400.275 ;
		RECT	0.255 247.485 0.57 247.635 ;
		RECT	0.255 403.005 0.57 403.155 ;
		RECT	0.255 405.885 0.57 406.035 ;
		RECT	0.255 408.765 0.57 408.915 ;
		RECT	0.255 411.645 0.57 411.795 ;
		RECT	0.255 250.365 0.57 250.515 ;
		RECT	0.255 253.245 0.57 253.395 ;
		RECT	0.255 256.125 0.57 256.275 ;
		RECT	15.63 187.305 16.17 187.415 ;
		RECT	15.63 185.175 16.17 186.575 ;
		RECT	16.17 187.305 16.71 187.415 ;
		RECT	16.17 185.175 16.71 186.575 ;
		RECT	16.71 187.305 17.25 187.415 ;
		RECT	16.71 185.175 17.25 186.575 ;
		RECT	15.09 187.305 15.63 187.415 ;
		RECT	15.09 185.175 15.63 186.575 ;
		RECT	14.49 187.305 15.09 187.415 ;
		RECT	14.49 185.175 15.09 186.575 ;
		RECT	17.25 187.305 17.79 187.415 ;
		RECT	17.25 185.175 17.79 186.575 ;
		RECT	17.79 187.305 18.33 187.415 ;
		RECT	17.79 185.175 18.33 186.575 ;
		RECT	18.33 187.305 18.87 187.415 ;
		RECT	18.33 185.175 18.87 186.575 ;
		RECT	19.41 187.305 20.01 187.415 ;
		RECT	19.41 185.175 20.01 186.575 ;
		RECT	18.87 187.305 19.41 187.415 ;
		RECT	18.87 185.175 19.41 186.575 ;
		RECT	15.09 227.445 15.63 227.555 ;
		RECT	15.09 228.285 15.63 229.685 ;
		RECT	14.49 227.445 15.09 227.555 ;
		RECT	14.49 228.285 15.09 229.685 ;
		RECT	15.63 227.445 16.17 227.555 ;
		RECT	15.63 228.285 16.17 229.685 ;
		RECT	16.17 227.445 16.71 227.555 ;
		RECT	16.17 228.285 16.71 229.685 ;
		RECT	16.71 227.445 17.25 227.555 ;
		RECT	16.71 228.285 17.25 229.685 ;
		RECT	17.25 227.445 17.79 227.555 ;
		RECT	17.25 228.285 17.79 229.685 ;
		RECT	17.79 227.445 18.33 227.555 ;
		RECT	17.79 228.285 18.33 229.685 ;
		RECT	18.33 227.445 18.87 227.555 ;
		RECT	18.33 228.285 18.87 229.685 ;
		RECT	19.41 227.445 20.01 227.555 ;
		RECT	19.41 228.285 20.01 229.685 ;
		RECT	18.87 227.445 19.41 227.555 ;
		RECT	18.87 228.285 19.41 229.685 ;
		RECT	20.01 185.175 21.165 186.575 ;
		RECT	20.01 187.305 21.165 187.415 ;
		RECT	20.97 187.415 21.165 187.835 ;
		RECT	20.01 187.55 20.87 187.74 ;
		RECT	20.01 188.225 21.165 188.325 ;
		RECT	20.01 189.205 21.165 189.31 ;
		RECT	20.97 189.31 21.165 189.655 ;
		RECT	20.01 189.41 20.87 189.6 ;
		RECT	20.97 189.835 21.165 190.175 ;
		RECT	20.01 189.885 20.87 190.075 ;
		RECT	20.92 190.175 21.165 190.33 ;
		RECT	20.01 190.18 20.86 190.33 ;
		RECT	20.01 190.72 21.165 190.785 ;
		RECT	20.01 191.175 21.165 191.28 ;
		RECT	20.01 191.67 21.165 191.77 ;
		RECT	20.41 192.16 21.165 192.26 ;
		RECT	20.01 192.65 21.165 192.755 ;
		RECT	20.79 192.755 21.165 193.145 ;
		RECT	20.01 193.145 21.165 193.245 ;
		RECT	20.01 193.635 21.165 193.74 ;
		RECT	20.97 193.74 21.165 194.13 ;
		RECT	20.01 193.84 20.87 194.03 ;
		RECT	20.01 194.13 21.165 194.23 ;
		RECT	20.01 194.62 21.165 194.725 ;
		RECT	20.01 195.115 21.165 195.215 ;
		RECT	20.01 195.605 21.165 195.705 ;
		RECT	20.01 196.095 21.165 196.2 ;
		RECT	20.01 196.59 21.165 196.69 ;
		RECT	20.01 197.08 21.165 197.18 ;
		RECT	20.01 197.57 21.165 197.675 ;
		RECT	20.97 197.675 21.165 198.065 ;
		RECT	20.01 197.775 20.87 197.965 ;
		RECT	20.01 198.065 21.165 198.165 ;
		RECT	20.01 198.555 21.165 198.66 ;
		RECT	20.01 199.05 21.165 199.15 ;
		RECT	20.01 199.54 21.165 199.63 ;
		RECT	20.01 200.04 21.165 200.135 ;
		RECT	20.01 200.525 21.165 200.625 ;
		RECT	20.01 201.015 21.165 201.12 ;
		RECT	20.01 201.51 21.165 201.6 ;
		RECT	20.97 201.6 21.165 202.01 ;
		RECT	20.01 201.7 20.87 201.91 ;
		RECT	20.01 202.01 21.165 202.105 ;
		RECT	20.97 202.105 21.165 202.495 ;
		RECT	20.01 202.495 21.165 202.6 ;
		RECT	20.01 202.99 21.165 203.085 ;
		RECT	20.01 203.475 21.165 203.58 ;
		RECT	20.01 203.97 21.165 204.055 ;
		RECT	20.97 204.055 21.165 205.055 ;
		RECT	20.01 204.455 20.87 204.665 ;
		RECT	20.01 204.78 20.86 204.97 ;
		RECT	20.97 205.59 21.165 205.895 ;
		RECT	20.01 205.645 20.87 205.835 ;
		RECT	20.01 206.43 21.165 206.53 ;
		RECT	20.01 206.92 21.165 207.02 ;
		RECT	20.01 207.41 21.165 207.515 ;
		RECT	20.01 207.905 21.165 208.005 ;
		RECT	20.01 208.395 21.165 208.5 ;
		RECT	20.97 209.035 21.165 209.335 ;
		RECT	20.01 209.09 20.87 209.28 ;
		RECT	20.97 209.87 21.165 210.87 ;
		RECT	20.01 209.895 20.87 210.085 ;
		RECT	20.01 210.23 20.87 210.44 ;
		RECT	20.01 210.87 21.165 210.955 ;
		RECT	20.01 211.345 21.165 211.45 ;
		RECT	20.01 211.84 21.165 211.945 ;
		RECT	20.01 212.335 21.165 212.425 ;
		RECT	20.97 212.425 21.165 212.835 ;
		RECT	20.01 212.835 21.165 212.915 ;
		RECT	20.97 212.915 21.165 213.325 ;
		RECT	20.01 213.015 20.87 213.225 ;
		RECT	20.01 213.325 21.165 213.42 ;
		RECT	20.01 213.81 21.165 213.91 ;
		RECT	20.01 214.3 21.165 214.405 ;
		RECT	20.01 214.795 21.165 214.885 ;
		RECT	20.01 215.295 21.165 215.385 ;
		RECT	20.01 215.775 21.165 215.88 ;
		RECT	20.01 216.27 21.165 216.37 ;
		RECT	20.01 216.76 21.165 216.865 ;
		RECT	20.97 216.865 21.165 217.255 ;
		RECT	20.01 216.965 20.87 217.155 ;
		RECT	20.01 217.255 21.165 217.355 ;
		RECT	20.01 217.745 21.165 217.845 ;
		RECT	20.01 218.235 21.165 218.34 ;
		RECT	20.01 218.73 21.165 218.83 ;
		RECT	20.01 219.22 21.165 219.325 ;
		RECT	20.01 219.715 21.165 219.815 ;
		RECT	20.01 220.205 21.165 220.305 ;
		RECT	20.41 220.695 21.165 220.79 ;
		RECT	20.97 220.79 21.165 221.2 ;
		RECT	20.01 220.89 20.87 221.1 ;
		RECT	20.01 221.2 21.165 221.29 ;
		RECT	20.01 221.68 21.165 221.775 ;
		RECT	20.79 221.775 21.165 222.185 ;
		RECT	20.74 222.185 21.165 222.275 ;
		RECT	20.74 222.665 21.165 222.755 ;
		RECT	20.01 223.165 21.165 223.225 ;
		RECT	20.01 223.615 21.165 223.75 ;
		RECT	20.01 224.14 21.165 224.21 ;
		RECT	20.97 224.6 21.165 225.09 ;
		RECT	20.01 224.6 20.87 224.75 ;
		RECT	20.01 224.85 20.87 225.04 ;
		RECT	20.97 225.27 21.165 225.615 ;
		RECT	20.01 225.325 20.87 225.515 ;
		RECT	20.01 225.615 21.165 225.72 ;
		RECT	20.01 226.6 21.165 226.705 ;
		RECT	20.97 227.095 21.165 227.445 ;
		RECT	20.01 227.105 20.87 227.315 ;
		RECT	20.01 227.445 21.165 227.555 ;
		RECT	20.01 228.285 21.165 229.685 ;
		RECT	14.49 187.55 19.41 187.74 ;
		RECT	14.49 188.225 19.41 188.325 ;
		RECT	14.49 189.205 19.41 189.31 ;
		RECT	14.49 189.41 19.41 189.6 ;
		RECT	14.49 189.885 19.41 190.075 ;
		RECT	14.59 190.18 19.41 190.33 ;
		RECT	14.49 190.72 19.41 190.785 ;
		RECT	14.49 191.175 19.41 191.28 ;
		RECT	14.49 191.67 19.41 191.77 ;
		RECT	14.49 192.65 19.41 192.755 ;
		RECT	14.49 193.145 19.41 193.245 ;
		RECT	14.49 193.635 19.41 193.74 ;
		RECT	14.49 193.84 19.41 194.03 ;
		RECT	14.49 194.13 19.41 194.23 ;
		RECT	14.49 194.62 19.41 194.725 ;
		RECT	14.49 195.115 19.41 195.215 ;
		RECT	14.49 195.605 19.41 195.705 ;
		RECT	14.49 196.095 19.41 196.2 ;
		RECT	14.49 196.59 19.41 196.69 ;
		RECT	14.49 197.08 19.41 197.18 ;
		RECT	14.49 197.57 19.41 197.675 ;
		RECT	14.49 197.775 19.41 197.965 ;
		RECT	14.49 198.065 19.41 198.165 ;
		RECT	14.49 198.555 19.41 198.66 ;
		RECT	14.49 199.05 19.41 199.15 ;
		RECT	14.49 199.54 19.41 199.63 ;
		RECT	14.49 200.04 19.41 200.135 ;
		RECT	14.49 200.525 19.41 200.625 ;
		RECT	14.49 201.015 19.41 201.12 ;
		RECT	14.49 201.51 19.41 201.6 ;
		RECT	14.49 201.7 19.41 201.91 ;
		RECT	14.49 202.01 19.41 202.105 ;
		RECT	14.49 202.495 19.41 202.6 ;
		RECT	14.49 202.99 19.41 203.085 ;
		RECT	14.49 203.475 19.41 203.58 ;
		RECT	14.49 203.97 19.41 204.055 ;
		RECT	14.49 204.445 14.595 204.68 ;
		RECT	14.695 204.455 19.41 204.665 ;
		RECT	14.49 204.78 19.41 204.97 ;
		RECT	14.49 205.645 19.41 205.835 ;
		RECT	14.49 206.43 19.41 206.53 ;
		RECT	14.49 206.92 19.41 207.02 ;
		RECT	14.49 207.41 19.41 207.515 ;
		RECT	14.49 207.905 19.41 208.005 ;
		RECT	14.49 208.395 19.41 208.5 ;
		RECT	14.49 209.09 19.41 209.28 ;
		RECT	14.49 209.895 19.41 210.085 ;
		RECT	14.59 210.23 19.41 210.44 ;
		RECT	14.49 210.87 19.41 210.955 ;
		RECT	14.49 211.345 19.41 211.45 ;
		RECT	14.49 211.84 19.41 211.945 ;
		RECT	14.49 212.335 19.41 212.425 ;
		RECT	14.49 212.835 19.41 212.915 ;
		RECT	14.49 213.015 19.41 213.225 ;
		RECT	14.49 213.325 19.41 213.42 ;
		RECT	14.49 213.81 19.41 213.91 ;
		RECT	14.49 214.3 19.41 214.405 ;
		RECT	14.49 214.795 19.41 214.885 ;
		RECT	14.49 215.295 19.41 215.385 ;
		RECT	14.49 215.775 19.41 215.88 ;
		RECT	14.49 216.27 19.41 216.37 ;
		RECT	14.49 216.76 19.41 216.865 ;
		RECT	14.49 216.965 19.41 217.155 ;
		RECT	14.49 217.255 19.41 217.355 ;
		RECT	14.49 217.745 19.41 217.845 ;
		RECT	14.49 218.235 19.41 218.34 ;
		RECT	14.49 218.73 19.41 218.83 ;
		RECT	14.49 219.22 19.41 219.325 ;
		RECT	14.49 219.715 19.41 219.815 ;
		RECT	14.49 220.205 19.41 220.305 ;
		RECT	14.49 220.89 19.41 221.1 ;
		RECT	14.49 221.2 19.41 221.29 ;
		RECT	14.49 221.68 19.41 221.775 ;
		RECT	14.49 222.19 19.41 222.26 ;
		RECT	14.49 222.68 19.445 222.75 ;
		RECT	14.49 223.165 19.41 223.225 ;
		RECT	14.49 223.615 19.41 223.75 ;
		RECT	14.49 224.14 19.41 224.21 ;
		RECT	14.49 224.6 14.63 224.75 ;
		RECT	14.69 224.6 19.41 224.75 ;
		RECT	14.49 224.85 19.41 225.04 ;
		RECT	14.49 225.325 19.41 225.515 ;
		RECT	14.49 225.615 19.41 225.72 ;
		RECT	14.49 226.6 19.41 226.705 ;
		RECT	14.49 227.105 19.41 227.315 ;
		RECT	19.41 187.55 20.01 187.74 ;
		RECT	19.41 188.225 20.01 188.325 ;
		RECT	19.41 189.205 20.01 189.31 ;
		RECT	19.41 189.41 20.01 189.6 ;
		RECT	19.41 189.885 20.01 190.075 ;
		RECT	19.41 190.18 20.175 190.33 ;
		RECT	19.41 190.72 20.01 190.785 ;
		RECT	19.41 191.175 20.01 191.28 ;
		RECT	19.41 191.67 20.01 191.77 ;
		RECT	19.41 192.65 20.01 192.755 ;
		RECT	19.41 193.145 20.01 193.245 ;
		RECT	19.41 193.635 20.01 193.74 ;
		RECT	19.41 193.84 20.01 194.03 ;
		RECT	19.41 194.13 20.01 194.23 ;
		RECT	19.41 194.62 20.01 194.725 ;
		RECT	19.41 195.115 20.01 195.215 ;
		RECT	19.41 195.605 20.01 195.705 ;
		RECT	19.41 196.095 20.01 196.2 ;
		RECT	19.41 196.59 20.01 196.69 ;
		RECT	19.41 197.08 20.01 197.18 ;
		RECT	19.41 197.57 20.01 197.675 ;
		RECT	19.41 197.775 20.01 197.965 ;
		RECT	19.41 198.065 20.01 198.165 ;
		RECT	19.41 198.555 20.01 198.66 ;
		RECT	19.41 199.05 20.01 199.15 ;
		RECT	19.41 199.54 20.01 199.63 ;
		RECT	19.41 200.04 20.01 200.135 ;
		RECT	19.41 200.525 20.01 200.625 ;
		RECT	19.41 201.015 20.01 201.12 ;
		RECT	19.41 201.51 20.01 201.6 ;
		RECT	19.41 201.7 20.01 201.91 ;
		RECT	19.41 202.01 20.01 202.105 ;
		RECT	19.41 202.495 20.01 202.6 ;
		RECT	19.41 202.99 20.01 203.085 ;
		RECT	19.41 203.475 20.01 203.58 ;
		RECT	19.41 203.97 20.01 204.055 ;
		RECT	19.41 204.455 20.085 204.665 ;
		RECT	19.41 204.78 20.01 204.97 ;
		RECT	19.41 205.645 20.01 205.835 ;
		RECT	19.41 206.43 20.01 206.53 ;
		RECT	19.41 206.92 20.01 207.02 ;
		RECT	19.41 207.41 20.01 207.515 ;
		RECT	19.41 207.905 20.01 208.005 ;
		RECT	19.41 208.395 20.01 208.5 ;
		RECT	19.41 209.09 20.01 209.28 ;
		RECT	19.41 209.895 20.01 210.085 ;
		RECT	19.41 210.23 20.01 210.44 ;
		RECT	19.41 210.87 20.01 210.955 ;
		RECT	19.41 211.345 20.01 211.45 ;
		RECT	19.41 211.84 20.01 211.945 ;
		RECT	19.41 212.335 20.01 212.425 ;
		RECT	19.41 212.835 20.01 212.915 ;
		RECT	19.41 213.015 20.01 213.225 ;
		RECT	19.41 213.325 20.01 213.42 ;
		RECT	19.41 213.81 20.01 213.91 ;
		RECT	19.41 214.3 20.01 214.405 ;
		RECT	19.41 214.795 20.01 214.885 ;
		RECT	19.41 215.295 20.01 215.385 ;
		RECT	19.41 215.775 20.01 215.88 ;
		RECT	19.41 216.27 20.01 216.37 ;
		RECT	19.41 216.76 20.01 216.865 ;
		RECT	19.41 216.965 20.01 217.155 ;
		RECT	19.41 217.255 20.01 217.355 ;
		RECT	19.41 217.745 20.01 217.845 ;
		RECT	19.41 218.235 20.01 218.34 ;
		RECT	19.41 218.73 20.01 218.83 ;
		RECT	19.41 219.22 20.01 219.325 ;
		RECT	19.41 219.715 20.01 219.815 ;
		RECT	19.41 220.205 20.01 220.305 ;
		RECT	19.41 220.89 20.01 221.1 ;
		RECT	19.41 221.2 20.01 221.29 ;
		RECT	19.41 221.68 20.01 221.775 ;
		RECT	19.41 222.19 20.01 222.26 ;
		RECT	19.41 222.68 20.01 222.75 ;
		RECT	19.41 223.165 20.01 223.225 ;
		RECT	19.41 223.615 20.01 223.75 ;
		RECT	19.41 224.14 20.01 224.21 ;
		RECT	19.41 224.6 20.01 224.75 ;
		RECT	19.41 224.85 20.01 225.04 ;
		RECT	19.41 225.325 20.01 225.515 ;
		RECT	19.41 225.615 20.01 225.72 ;
		RECT	19.41 226.6 20.01 226.705 ;
		RECT	19.41 227.105 20.01 227.315 ;
		RECT	0.295 192.855 20.69 193.045 ;
		RECT	0.215 202.205 20.87 202.395 ;
		RECT	0.21 204.155 20.86 204.345 ;
		RECT	0.22 210.58 20.87 210.77 ;
		RECT	0.225 212.525 20.87 212.735 ;
		RECT	0.225 221.875 20.69 222.085 ;
		RECT	0.225 222.19 0.57 222.26 ;
		RECT	0.22 222.68 0.57 222.75 ;
		RECT	11.61 188.72 21.07 188.81 ;
		RECT	11.61 189.705 21.07 189.785 ;
		RECT	14.2 192.165 20.36 192.255 ;
		RECT	13.85 205.45 21.07 205.54 ;
		RECT	13.85 205.945 21.07 206.035 ;
		RECT	7.07 207.415 13.545 207.515 ;
		RECT	13.85 208.895 21.07 208.985 ;
		RECT	13.85 209.385 21.07 209.475 ;
		RECT	14.2 220.7 20.36 220.79 ;
		RECT	0.57 221.205 2.735 221.275 ;
		RECT	12.605 225.14 21.07 225.22 ;
		RECT	12.605 226.115 21.07 226.205 ;
		RECT	20.01 222.19 20.69 222.26 ;
		RECT	20.01 222.68 20.69 222.75 ;
		LAYER	VIA1 DESIGNRULEWIDTH 0.07 ;
		RECT	0 0 21.165 414.86 ;
		LAYER	VIA2 DESIGNRULEWIDTH 0.07 ;
		RECT	0 0 21.165 414.86 ;
		LAYER	VIA3 DESIGNRULEWIDTH 0.07 ;
		RECT	0.435 186.415 0.485 186.545 ;
		RECT	0.435 187.58 0.485 187.71 ;
		RECT	0.435 189.445 0.485 189.575 ;
		RECT	0.435 189.915 0.485 190.045 ;
		RECT	0.435 193.87 0.485 194 ;
		RECT	0.435 197.805 0.485 197.935 ;
		RECT	0.435 201.74 0.485 201.87 ;
		RECT	0.435 204.865 0.485 204.995 ;
		RECT	0.435 205.675 0.485 205.805 ;
		RECT	0.435 209.12 0.485 209.25 ;
		RECT	0.435 209.93 0.485 210.06 ;
		RECT	0.435 213.055 0.485 213.185 ;
		RECT	0.435 216.995 0.485 217.125 ;
		RECT	0.435 220.93 0.485 221.06 ;
		RECT	0.435 224.88 0.485 225.01 ;
		RECT	0.435 225.355 0.485 225.485 ;
		RECT	0.435 227.145 0.485 227.275 ;
		RECT	0.435 228.315 0.485 228.445 ;
		RECT	0.435 186.875 0.485 187.005 ;
		RECT	0.435 192.885 0.485 193.015 ;
		RECT	0.435 221.915 0.485 222.045 ;
		RECT	0.435 227.855 0.485 227.985 ;
		RECT	1.085 186.415 1.135 186.545 ;
		RECT	1.38 186.415 1.43 186.545 ;
		RECT	1.86 186.415 1.91 186.545 ;
		RECT	2.01 186.415 2.06 186.545 ;
		RECT	3.25 186.415 3.3 186.545 ;
		RECT	3.515 186.415 3.565 186.545 ;
		RECT	4.51 186.415 4.56 186.545 ;
		RECT	5.035 186.415 5.085 186.545 ;
		RECT	6.22 186.415 6.27 186.545 ;
		RECT	7.5 186.415 7.55 186.545 ;
		RECT	9.315 186.415 9.365 186.545 ;
		RECT	9.72 186.415 9.77 186.545 ;
		RECT	11.025 186.415 11.075 186.545 ;
		RECT	0.62 186.645 0.67 186.775 ;
		RECT	3.65 186.645 3.7 186.775 ;
		RECT	7.19 186.645 7.24 186.775 ;
		RECT	14.14 186.645 14.19 186.775 ;
		RECT	2.18 186.875 2.23 187.005 ;
		RECT	8.56 186.875 8.61 187.005 ;
		RECT	10.27 186.875 10.32 187.005 ;
		RECT	13.8 187.105 13.85 187.235 ;
		RECT	1.045 187.555 1.175 187.605 ;
		RECT	1.34 187.555 1.47 187.605 ;
		RECT	4.47 187.555 4.6 187.605 ;
		RECT	9.275 187.555 9.405 187.605 ;
		RECT	1.86 187.58 1.91 187.71 ;
		RECT	2.01 187.58 2.06 187.71 ;
		RECT	3.25 187.58 3.3 187.71 ;
		RECT	3.515 187.58 3.565 187.71 ;
		RECT	5.035 187.58 5.085 187.71 ;
		RECT	6.22 187.58 6.27 187.71 ;
		RECT	7.5 187.58 7.55 187.71 ;
		RECT	9.72 187.58 9.77 187.71 ;
		RECT	11.025 187.58 11.075 187.71 ;
		RECT	1.045 187.685 1.175 187.735 ;
		RECT	1.34 187.685 1.47 187.735 ;
		RECT	4.47 187.685 4.6 187.735 ;
		RECT	9.275 187.685 9.405 187.735 ;
		RECT	3.02 187.94 3.15 187.99 ;
		RECT	1.57 187.965 1.62 188.095 ;
		RECT	4.87 187.965 4.92 188.095 ;
		RECT	5.9 187.965 5.95 188.095 ;
		RECT	8.955 187.965 9.005 188.095 ;
		RECT	12.79 187.965 12.84 188.095 ;
		RECT	14.33 187.965 14.38 188.095 ;
		RECT	3.02 188.07 3.15 188.12 ;
		RECT	3.8 188.43 3.93 188.48 ;
		RECT	5.635 188.43 5.765 188.48 ;
		RECT	8.31 188.43 8.44 188.48 ;
		RECT	8.73 188.43 8.86 188.48 ;
		RECT	0.9 188.455 0.95 188.585 ;
		RECT	2.485 188.455 2.535 188.585 ;
		RECT	2.615 188.455 2.665 188.585 ;
		RECT	6.065 188.455 6.115 188.585 ;
		RECT	6.725 188.455 6.775 188.585 ;
		RECT	11.555 188.455 11.865 188.585 ;
		RECT	12.52 188.455 12.57 188.585 ;
		RECT	14.005 188.455 14.055 188.585 ;
		RECT	3.8 188.56 3.93 188.61 ;
		RECT	5.635 188.56 5.765 188.61 ;
		RECT	8.31 188.56 8.44 188.61 ;
		RECT	8.73 188.56 8.86 188.61 ;
		RECT	11.685 188.74 11.735 188.79 ;
		RECT	12.655 188.74 12.705 188.79 ;
		RECT	3.02 188.92 3.15 188.97 ;
		RECT	1.57 188.945 1.62 189.075 ;
		RECT	4.87 188.945 4.92 189.075 ;
		RECT	5.9 188.945 5.95 189.075 ;
		RECT	8.955 188.945 9.005 189.075 ;
		RECT	12.79 188.945 12.84 189.075 ;
		RECT	14.335 188.945 14.385 189.075 ;
		RECT	3.02 189.05 3.15 189.1 ;
		RECT	1.045 189.42 1.175 189.47 ;
		RECT	1.34 189.42 1.47 189.47 ;
		RECT	4.47 189.42 4.6 189.47 ;
		RECT	9.275 189.42 9.405 189.47 ;
		RECT	13.675 189.44 13.725 189.57 ;
		RECT	1.86 189.445 1.91 189.575 ;
		RECT	2.01 189.445 2.06 189.575 ;
		RECT	3.25 189.445 3.3 189.575 ;
		RECT	3.515 189.445 3.565 189.575 ;
		RECT	5.035 189.445 5.085 189.575 ;
		RECT	6.22 189.445 6.27 189.575 ;
		RECT	7.5 189.445 7.55 189.575 ;
		RECT	9.72 189.445 9.77 189.575 ;
		RECT	11.025 189.445 11.075 189.575 ;
		RECT	1.045 189.55 1.175 189.6 ;
		RECT	1.34 189.55 1.47 189.6 ;
		RECT	4.47 189.55 4.6 189.6 ;
		RECT	9.275 189.55 9.405 189.6 ;
		RECT	11.685 189.72 11.735 189.77 ;
		RECT	12.655 189.72 12.705 189.77 ;
		RECT	1.045 189.89 1.175 189.94 ;
		RECT	1.34 189.89 1.47 189.94 ;
		RECT	4.47 189.89 4.6 189.94 ;
		RECT	9.275 189.89 9.405 189.94 ;
		RECT	1.86 189.915 1.91 190.045 ;
		RECT	2.01 189.915 2.06 190.045 ;
		RECT	3.25 189.915 3.3 190.045 ;
		RECT	3.515 189.915 3.565 190.045 ;
		RECT	5.035 189.915 5.085 190.045 ;
		RECT	6.22 189.915 6.27 190.045 ;
		RECT	7.5 189.915 7.55 190.045 ;
		RECT	9.72 189.915 9.77 190.045 ;
		RECT	11.025 189.915 11.075 190.045 ;
		RECT	1.045 190.02 1.175 190.07 ;
		RECT	1.34 190.02 1.47 190.07 ;
		RECT	4.47 190.02 4.6 190.07 ;
		RECT	9.275 190.02 9.405 190.07 ;
		RECT	3.8 190.435 3.93 190.485 ;
		RECT	5.635 190.435 5.765 190.485 ;
		RECT	8.31 190.435 8.44 190.485 ;
		RECT	8.73 190.435 8.86 190.485 ;
		RECT	0.9 190.46 0.95 190.59 ;
		RECT	2.485 190.46 2.535 190.59 ;
		RECT	2.615 190.46 2.665 190.59 ;
		RECT	6.065 190.46 6.115 190.59 ;
		RECT	6.725 190.46 6.775 190.59 ;
		RECT	11.555 190.46 11.865 190.59 ;
		RECT	12.52 190.46 12.57 190.59 ;
		RECT	14.005 190.46 14.055 190.59 ;
		RECT	3.8 190.565 3.93 190.615 ;
		RECT	5.635 190.565 5.765 190.615 ;
		RECT	8.31 190.565 8.44 190.615 ;
		RECT	8.73 190.565 8.86 190.615 ;
		RECT	3.02 190.89 3.15 190.94 ;
		RECT	1.57 190.915 1.62 191.045 ;
		RECT	4.87 190.915 4.92 191.045 ;
		RECT	5.9 190.915 5.95 191.045 ;
		RECT	8.955 190.915 9.005 191.045 ;
		RECT	12.79 190.915 12.84 191.045 ;
		RECT	14.335 190.915 14.385 191.045 ;
		RECT	3.02 191.02 3.15 191.07 ;
		RECT	4.035 191.41 4.085 191.54 ;
		RECT	6.495 191.41 6.545 191.54 ;
		RECT	11.685 191.41 11.735 191.54 ;
		RECT	12.655 191.41 12.705 191.54 ;
		RECT	3.02 191.875 3.15 191.925 ;
		RECT	1.57 191.9 1.62 192.03 ;
		RECT	4.87 191.9 4.92 192.03 ;
		RECT	5.9 191.9 5.95 192.03 ;
		RECT	8.955 191.9 9.005 192.03 ;
		RECT	12.79 191.9 12.84 192.03 ;
		RECT	14.335 191.9 14.385 192.03 ;
		RECT	3.02 192.005 3.15 192.055 ;
		RECT	14.29 192.185 14.42 192.235 ;
		RECT	4.035 192.39 4.085 192.52 ;
		RECT	6.495 192.39 6.545 192.52 ;
		RECT	2.18 192.885 2.23 193.015 ;
		RECT	8.56 192.885 8.61 193.015 ;
		RECT	10.27 192.885 10.32 193.015 ;
		RECT	3.8 193.35 3.93 193.4 ;
		RECT	5.635 193.35 5.765 193.4 ;
		RECT	8.31 193.35 8.44 193.4 ;
		RECT	8.73 193.35 8.86 193.4 ;
		RECT	0.9 193.375 0.95 193.505 ;
		RECT	2.485 193.375 2.535 193.505 ;
		RECT	2.615 193.375 2.665 193.505 ;
		RECT	6.065 193.375 6.115 193.505 ;
		RECT	6.725 193.375 6.775 193.505 ;
		RECT	11.555 193.375 11.865 193.505 ;
		RECT	12.52 193.375 12.57 193.505 ;
		RECT	14.005 193.375 14.055 193.505 ;
		RECT	3.8 193.48 3.93 193.53 ;
		RECT	5.635 193.48 5.765 193.53 ;
		RECT	8.31 193.48 8.44 193.53 ;
		RECT	8.73 193.48 8.86 193.53 ;
		RECT	1.045 193.845 1.175 193.895 ;
		RECT	1.34 193.845 1.47 193.895 ;
		RECT	4.47 193.845 4.6 193.895 ;
		RECT	1.86 193.87 1.91 194 ;
		RECT	2.01 193.87 2.06 194 ;
		RECT	2.32 193.87 2.37 194 ;
		RECT	3.25 193.87 3.3 194 ;
		RECT	3.515 193.87 3.565 194 ;
		RECT	5.035 193.87 5.085 194 ;
		RECT	6.22 193.87 6.27 194 ;
		RECT	7.5 193.87 7.55 194 ;
		RECT	9.72 193.87 9.77 194 ;
		RECT	11.025 193.87 11.075 194 ;
		RECT	1.045 193.975 1.175 194.025 ;
		RECT	1.34 193.975 1.47 194.025 ;
		RECT	4.47 193.975 4.6 194.025 ;
		RECT	3.8 194.335 3.93 194.385 ;
		RECT	5.635 194.335 5.765 194.385 ;
		RECT	8.31 194.335 8.44 194.385 ;
		RECT	8.73 194.335 8.86 194.385 ;
		RECT	0.9 194.36 0.95 194.49 ;
		RECT	2.485 194.36 2.535 194.49 ;
		RECT	2.615 194.36 2.665 194.49 ;
		RECT	6.065 194.36 6.115 194.49 ;
		RECT	6.725 194.36 6.775 194.49 ;
		RECT	11.555 194.36 11.865 194.49 ;
		RECT	12.52 194.36 12.57 194.49 ;
		RECT	14.005 194.36 14.055 194.49 ;
		RECT	3.8 194.465 3.93 194.515 ;
		RECT	5.635 194.465 5.765 194.515 ;
		RECT	8.31 194.465 8.44 194.515 ;
		RECT	8.73 194.465 8.86 194.515 ;
		RECT	3.02 194.83 3.15 194.88 ;
		RECT	1.57 194.855 1.62 194.985 ;
		RECT	4.87 194.855 4.92 194.985 ;
		RECT	5.9 194.855 5.95 194.985 ;
		RECT	9.195 194.855 9.245 194.985 ;
		RECT	10.27 194.855 10.32 194.985 ;
		RECT	12.79 194.855 12.84 194.985 ;
		RECT	14.335 194.855 14.385 194.985 ;
		RECT	3.02 194.96 3.15 195.01 ;
		RECT	4.035 195.345 4.085 195.475 ;
		RECT	3.02 195.81 3.15 195.86 ;
		RECT	1.57 195.835 1.62 195.965 ;
		RECT	4.87 195.835 4.92 195.965 ;
		RECT	5.9 195.835 5.95 195.965 ;
		RECT	9.195 195.835 9.245 195.965 ;
		RECT	9.43 195.835 9.48 195.965 ;
		RECT	10.27 195.835 10.32 195.965 ;
		RECT	12.79 195.835 12.84 195.965 ;
		RECT	14.335 195.835 14.385 195.965 ;
		RECT	3.02 195.94 3.15 195.99 ;
		RECT	0.9 196.305 14.055 196.485 ;
		RECT	3.02 196.795 3.15 196.845 ;
		RECT	1.57 196.82 1.62 196.95 ;
		RECT	4.87 196.82 4.92 196.95 ;
		RECT	5.9 196.82 5.95 196.95 ;
		RECT	9.43 196.82 9.48 196.95 ;
		RECT	10.27 196.82 10.32 196.95 ;
		RECT	12.79 196.82 12.84 196.95 ;
		RECT	14.33 196.82 14.38 196.95 ;
		RECT	3.02 196.925 3.15 196.975 ;
		RECT	3.8 197.285 3.93 197.335 ;
		RECT	5.635 197.285 5.765 197.335 ;
		RECT	8.31 197.285 8.44 197.335 ;
		RECT	8.73 197.285 8.86 197.335 ;
		RECT	0.9 197.31 0.95 197.44 ;
		RECT	2.485 197.31 2.535 197.44 ;
		RECT	2.615 197.31 2.665 197.44 ;
		RECT	6.065 197.31 6.115 197.44 ;
		RECT	6.725 197.31 6.775 197.44 ;
		RECT	11.555 197.31 11.865 197.44 ;
		RECT	12.52 197.31 12.57 197.44 ;
		RECT	14.005 197.31 14.055 197.44 ;
		RECT	3.8 197.415 3.93 197.465 ;
		RECT	5.635 197.415 5.765 197.465 ;
		RECT	8.31 197.415 8.44 197.465 ;
		RECT	8.73 197.415 8.86 197.465 ;
		RECT	1.045 197.78 1.175 197.83 ;
		RECT	1.34 197.78 1.47 197.83 ;
		RECT	4.47 197.78 4.6 197.83 ;
		RECT	1.86 197.805 1.91 197.935 ;
		RECT	2.01 197.805 2.06 197.935 ;
		RECT	2.32 197.805 2.37 197.935 ;
		RECT	3.25 197.805 3.3 197.935 ;
		RECT	3.515 197.805 3.565 197.935 ;
		RECT	5.035 197.805 5.085 197.935 ;
		RECT	6.22 197.805 6.27 197.935 ;
		RECT	7.5 197.805 7.55 197.935 ;
		RECT	9.72 197.805 9.77 197.935 ;
		RECT	11.025 197.805 11.075 197.935 ;
		RECT	1.045 197.91 1.175 197.96 ;
		RECT	1.34 197.91 1.47 197.96 ;
		RECT	4.47 197.91 4.6 197.96 ;
		RECT	3.8 198.27 3.93 198.32 ;
		RECT	5.635 198.27 5.765 198.32 ;
		RECT	8.31 198.27 8.44 198.32 ;
		RECT	8.73 198.27 8.86 198.32 ;
		RECT	0.9 198.295 0.95 198.425 ;
		RECT	2.485 198.295 2.535 198.425 ;
		RECT	2.615 198.295 2.665 198.425 ;
		RECT	6.065 198.295 6.115 198.425 ;
		RECT	6.725 198.295 6.775 198.425 ;
		RECT	11.555 198.295 11.865 198.425 ;
		RECT	12.52 198.295 12.57 198.425 ;
		RECT	14.005 198.295 14.055 198.425 ;
		RECT	3.8 198.4 3.93 198.45 ;
		RECT	5.635 198.4 5.765 198.45 ;
		RECT	8.31 198.4 8.44 198.45 ;
		RECT	8.73 198.4 8.86 198.45 ;
		RECT	3.02 198.765 3.15 198.815 ;
		RECT	1.57 198.79 1.62 198.92 ;
		RECT	4.87 198.79 4.92 198.92 ;
		RECT	5.9 198.79 5.95 198.92 ;
		RECT	6.375 198.79 6.425 198.92 ;
		RECT	10.27 198.79 10.32 198.92 ;
		RECT	12.65 198.79 12.84 198.92 ;
		RECT	14.33 198.79 14.38 198.92 ;
		RECT	3.02 198.895 3.15 198.945 ;
		RECT	4.035 199.28 4.085 199.41 ;
		RECT	6.835 199.565 6.885 199.615 ;
		RECT	3.02 199.745 3.15 199.795 ;
		RECT	1.57 199.77 1.62 199.9 ;
		RECT	4.87 199.77 4.92 199.9 ;
		RECT	5.9 199.77 5.95 199.9 ;
		RECT	6.375 199.77 6.425 199.9 ;
		RECT	7.015 199.77 7.065 199.9 ;
		RECT	10.27 199.77 10.32 199.9 ;
		RECT	12.79 199.77 12.84 199.9 ;
		RECT	14.33 199.77 14.38 199.9 ;
		RECT	3.02 199.875 3.15 199.925 ;
		RECT	4.035 200.265 4.085 200.395 ;
		RECT	3.02 200.73 3.15 200.78 ;
		RECT	1.57 200.755 1.62 200.885 ;
		RECT	4.87 200.755 4.92 200.885 ;
		RECT	5.9 200.755 5.95 200.885 ;
		RECT	6.375 200.755 6.425 200.885 ;
		RECT	7.015 200.755 7.065 200.885 ;
		RECT	10.27 200.755 10.32 200.885 ;
		RECT	12.79 200.755 12.84 200.885 ;
		RECT	14.33 200.755 14.38 200.885 ;
		RECT	3.02 200.86 3.15 200.91 ;
		RECT	0.9 201.25 0.95 201.38 ;
		RECT	2.485 201.25 2.535 201.38 ;
		RECT	2.615 201.25 2.665 201.38 ;
		RECT	6.065 201.25 6.115 201.38 ;
		RECT	6.675 201.25 6.725 201.38 ;
		RECT	11.555 201.25 11.865 201.38 ;
		RECT	12.52 201.25 12.57 201.38 ;
		RECT	14.005 201.25 14.055 201.38 ;
		RECT	3.8 201.29 3.93 201.34 ;
		RECT	5.635 201.29 5.765 201.34 ;
		RECT	8.31 201.29 8.44 201.34 ;
		RECT	8.73 201.29 8.86 201.34 ;
		RECT	9.315 201.535 9.445 201.585 ;
		RECT	1.045 201.715 1.175 201.765 ;
		RECT	1.34 201.715 1.47 201.765 ;
		RECT	4.47 201.715 4.6 201.765 ;
		RECT	1.86 201.74 1.91 201.87 ;
		RECT	2.01 201.74 2.06 201.87 ;
		RECT	2.32 201.74 2.37 201.87 ;
		RECT	3.25 201.74 3.3 201.87 ;
		RECT	3.515 201.74 3.565 201.87 ;
		RECT	5.035 201.74 5.085 201.87 ;
		RECT	6.22 201.74 6.27 201.87 ;
		RECT	7.5 201.74 7.55 201.87 ;
		RECT	9.72 201.74 9.77 201.87 ;
		RECT	11.025 201.74 11.075 201.87 ;
		RECT	1.045 201.845 1.175 201.895 ;
		RECT	1.34 201.845 1.47 201.895 ;
		RECT	4.47 201.845 4.6 201.895 ;
		RECT	0.62 202.235 0.67 202.365 ;
		RECT	3.65 202.235 3.7 202.365 ;
		RECT	7.19 202.235 7.24 202.365 ;
		RECT	14.14 202.235 14.19 202.365 ;
		RECT	3.02 202.705 3.15 202.755 ;
		RECT	1.57 202.73 1.62 202.86 ;
		RECT	4.87 202.73 4.92 202.86 ;
		RECT	5.9 202.73 5.95 202.86 ;
		RECT	6.375 202.73 6.425 202.86 ;
		RECT	7.015 202.73 7.065 202.86 ;
		RECT	10.27 202.73 10.32 202.86 ;
		RECT	12.79 202.73 12.84 202.86 ;
		RECT	14.335 202.73 14.385 202.86 ;
		RECT	3.02 202.835 3.15 202.885 ;
		RECT	4.035 203.215 4.085 203.345 ;
		RECT	11.685 203.215 11.735 203.345 ;
		RECT	13.9 203.215 13.95 203.345 ;
		RECT	3.02 203.685 3.15 203.735 ;
		RECT	1.57 203.71 1.62 203.84 ;
		RECT	4.87 203.71 4.92 203.84 ;
		RECT	5.9 203.71 5.95 203.84 ;
		RECT	6.375 203.71 6.425 203.84 ;
		RECT	7.015 203.71 7.065 203.84 ;
		RECT	10.27 203.71 10.32 203.84 ;
		RECT	12.79 203.71 12.84 203.84 ;
		RECT	14.335 203.71 14.385 203.84 ;
		RECT	3.02 203.815 3.15 203.865 ;
		RECT	13.8 204.185 13.85 204.315 ;
		RECT	13.675 204.81 13.725 204.94 ;
		RECT	1.085 204.865 1.135 204.995 ;
		RECT	1.38 204.865 1.43 204.995 ;
		RECT	1.86 204.865 1.91 204.995 ;
		RECT	2.01 204.865 2.06 204.995 ;
		RECT	2.32 204.865 2.37 204.995 ;
		RECT	3.25 204.865 3.3 204.995 ;
		RECT	3.515 204.865 3.565 204.995 ;
		RECT	4.51 204.865 4.56 204.995 ;
		RECT	5.035 204.865 5.085 204.995 ;
		RECT	6.22 204.865 6.27 204.995 ;
		RECT	7.5 204.865 7.55 204.995 ;
		RECT	9.72 204.865 9.77 204.995 ;
		RECT	11.025 204.865 11.075 204.995 ;
		RECT	3.8 205.16 3.93 205.21 ;
		RECT	5.635 205.16 5.765 205.21 ;
		RECT	8.31 205.16 8.44 205.21 ;
		RECT	8.73 205.16 8.86 205.21 ;
		RECT	0.9 205.185 0.95 205.315 ;
		RECT	2.485 205.185 2.535 205.315 ;
		RECT	2.615 205.185 2.665 205.315 ;
		RECT	6.065 205.185 6.115 205.315 ;
		RECT	6.675 205.185 6.725 205.315 ;
		RECT	11.555 205.185 11.865 205.315 ;
		RECT	12.52 205.185 12.57 205.315 ;
		RECT	14.005 205.185 14.055 205.315 ;
		RECT	3.8 205.29 3.93 205.34 ;
		RECT	5.635 205.29 5.765 205.34 ;
		RECT	8.31 205.29 8.44 205.34 ;
		RECT	8.73 205.29 8.86 205.34 ;
		RECT	13.9 205.47 13.95 205.52 ;
		RECT	1.045 205.65 1.175 205.7 ;
		RECT	1.34 205.65 1.47 205.7 ;
		RECT	4.47 205.65 4.6 205.7 ;
		RECT	1.86 205.675 1.91 205.805 ;
		RECT	2.01 205.675 2.06 205.805 ;
		RECT	2.32 205.675 2.37 205.805 ;
		RECT	3.25 205.675 3.3 205.805 ;
		RECT	3.515 205.675 3.565 205.805 ;
		RECT	5.035 205.675 5.085 205.805 ;
		RECT	6.22 205.675 6.27 205.805 ;
		RECT	7.5 205.675 7.55 205.805 ;
		RECT	9.72 205.675 9.77 205.805 ;
		RECT	11.025 205.675 11.075 205.805 ;
		RECT	1.045 205.78 1.175 205.83 ;
		RECT	1.34 205.78 1.47 205.83 ;
		RECT	4.47 205.78 4.6 205.83 ;
		RECT	13.9 205.965 13.95 206.015 ;
		RECT	3.8 206.145 3.93 206.195 ;
		RECT	5.635 206.145 5.765 206.195 ;
		RECT	8.31 206.145 8.44 206.195 ;
		RECT	8.73 206.145 8.86 206.195 ;
		RECT	0.9 206.17 0.95 206.3 ;
		RECT	2.485 206.17 2.535 206.3 ;
		RECT	2.615 206.17 2.665 206.3 ;
		RECT	6.065 206.17 6.115 206.3 ;
		RECT	6.675 206.17 6.725 206.3 ;
		RECT	10.12 206.17 10.17 206.3 ;
		RECT	11.555 206.17 11.865 206.3 ;
		RECT	12.52 206.17 12.57 206.3 ;
		RECT	14.005 206.17 14.055 206.3 ;
		RECT	3.8 206.275 3.93 206.325 ;
		RECT	5.635 206.275 5.765 206.325 ;
		RECT	8.31 206.275 8.44 206.325 ;
		RECT	8.73 206.275 8.86 206.325 ;
		RECT	3.02 206.635 3.15 206.685 ;
		RECT	1.57 206.66 1.62 206.79 ;
		RECT	4.87 206.66 4.92 206.79 ;
		RECT	5.9 206.66 5.95 206.79 ;
		RECT	6.375 206.66 6.425 206.79 ;
		RECT	7.015 206.66 7.065 206.79 ;
		RECT	9.11 206.66 9.16 206.79 ;
		RECT	10.27 206.66 10.32 206.79 ;
		RECT	12.79 206.66 12.84 206.79 ;
		RECT	14.335 206.66 14.385 206.79 ;
		RECT	3.02 206.765 3.15 206.815 ;
		RECT	4.035 207.15 4.085 207.28 ;
		RECT	13.9 207.15 13.95 207.28 ;
		RECT	7.19 207.44 7.24 207.49 ;
		RECT	12.655 207.44 12.705 207.49 ;
		RECT	4.035 207.645 4.085 207.775 ;
		RECT	13.9 207.645 13.95 207.775 ;
		RECT	3.02 208.11 3.15 208.16 ;
		RECT	1.57 208.135 1.62 208.265 ;
		RECT	4.87 208.135 4.92 208.265 ;
		RECT	5.9 208.135 5.95 208.265 ;
		RECT	6.375 208.135 6.425 208.265 ;
		RECT	7.015 208.135 7.065 208.265 ;
		RECT	9.11 208.135 9.16 208.265 ;
		RECT	10.27 208.135 10.32 208.265 ;
		RECT	12.79 208.135 12.84 208.265 ;
		RECT	14.335 208.135 14.385 208.265 ;
		RECT	3.02 208.24 3.15 208.29 ;
		RECT	3.8 208.605 3.93 208.655 ;
		RECT	4.22 208.605 4.35 208.655 ;
		RECT	5.635 208.605 5.765 208.655 ;
		RECT	8.31 208.605 8.44 208.655 ;
		RECT	8.73 208.605 8.86 208.655 ;
		RECT	0.9 208.63 0.95 208.76 ;
		RECT	2.485 208.63 2.535 208.76 ;
		RECT	2.615 208.63 2.665 208.76 ;
		RECT	6.065 208.63 6.115 208.76 ;
		RECT	6.675 208.63 6.725 208.76 ;
		RECT	10.12 208.63 10.17 208.76 ;
		RECT	11.555 208.63 11.865 208.76 ;
		RECT	12.52 208.63 12.57 208.76 ;
		RECT	14.005 208.63 14.055 208.76 ;
		RECT	3.8 208.735 3.93 208.785 ;
		RECT	4.22 208.735 4.35 208.785 ;
		RECT	5.635 208.735 5.765 208.785 ;
		RECT	8.31 208.735 8.44 208.785 ;
		RECT	8.73 208.735 8.86 208.785 ;
		RECT	13.9 208.915 13.95 208.965 ;
		RECT	1.045 209.095 1.175 209.145 ;
		RECT	1.34 209.095 1.47 209.145 ;
		RECT	4.47 209.095 4.6 209.145 ;
		RECT	1.86 209.12 1.91 209.25 ;
		RECT	2.01 209.12 2.06 209.25 ;
		RECT	2.32 209.12 2.37 209.25 ;
		RECT	3.25 209.12 3.3 209.25 ;
		RECT	3.515 209.12 3.565 209.25 ;
		RECT	5.035 209.12 5.085 209.25 ;
		RECT	6.22 209.12 6.27 209.25 ;
		RECT	7.5 209.12 7.55 209.25 ;
		RECT	9.72 209.12 9.77 209.25 ;
		RECT	11.025 209.12 11.075 209.25 ;
		RECT	1.045 209.225 1.175 209.275 ;
		RECT	1.34 209.225 1.47 209.275 ;
		RECT	4.47 209.225 4.6 209.275 ;
		RECT	13.9 209.405 13.95 209.455 ;
		RECT	0.9 209.585 14.055 209.765 ;
		RECT	13.675 209.925 13.725 210.055 ;
		RECT	1.085 209.93 1.135 210.06 ;
		RECT	1.38 209.93 1.43 210.06 ;
		RECT	1.86 209.93 1.91 210.06 ;
		RECT	2.01 209.93 2.06 210.06 ;
		RECT	2.32 209.93 2.37 210.06 ;
		RECT	3.25 209.93 3.3 210.06 ;
		RECT	3.515 209.93 3.565 210.06 ;
		RECT	4.51 209.93 4.56 210.06 ;
		RECT	5.035 209.93 5.085 210.06 ;
		RECT	6.22 209.93 6.27 210.06 ;
		RECT	7.5 209.93 7.55 210.06 ;
		RECT	9.72 209.93 9.77 210.06 ;
		RECT	11.025 209.93 11.075 210.06 ;
		RECT	13.8 210.61 13.85 210.74 ;
		RECT	3.02 211.06 3.15 211.11 ;
		RECT	1.57 211.085 1.62 211.215 ;
		RECT	4.87 211.085 4.92 211.215 ;
		RECT	6.375 211.085 6.425 211.215 ;
		RECT	7.015 211.085 7.065 211.215 ;
		RECT	10.27 211.085 10.32 211.215 ;
		RECT	12.79 211.085 12.84 211.215 ;
		RECT	14.33 211.085 14.38 211.215 ;
		RECT	3.02 211.19 3.15 211.24 ;
		RECT	4.035 211.58 4.085 211.71 ;
		RECT	12.655 211.58 12.705 211.71 ;
		RECT	13.9 211.58 13.95 211.71 ;
		RECT	3.02 212.05 3.15 212.1 ;
		RECT	1.57 212.075 1.62 212.205 ;
		RECT	4.87 212.075 4.92 212.205 ;
		RECT	6.375 212.075 6.425 212.205 ;
		RECT	7.015 212.075 7.065 212.205 ;
		RECT	10.27 212.075 10.32 212.205 ;
		RECT	12.79 212.075 12.84 212.205 ;
		RECT	14.33 212.075 14.38 212.205 ;
		RECT	3.02 212.18 3.15 212.23 ;
		RECT	0.62 212.565 0.67 212.695 ;
		RECT	3.65 212.565 3.7 212.695 ;
		RECT	7.19 212.565 7.24 212.695 ;
		RECT	14.14 212.565 14.19 212.695 ;
		RECT	6.85 212.85 6.9 212.9 ;
		RECT	1.045 213.03 1.175 213.08 ;
		RECT	1.34 213.03 1.47 213.08 ;
		RECT	4.47 213.03 4.6 213.08 ;
		RECT	1.86 213.055 1.91 213.185 ;
		RECT	2.01 213.055 2.06 213.185 ;
		RECT	2.32 213.055 2.37 213.185 ;
		RECT	3.25 213.055 3.3 213.185 ;
		RECT	3.515 213.055 3.565 213.185 ;
		RECT	5.035 213.055 5.085 213.185 ;
		RECT	6.22 213.055 6.27 213.185 ;
		RECT	7.5 213.055 7.55 213.185 ;
		RECT	9.72 213.055 9.77 213.185 ;
		RECT	11.025 213.055 11.075 213.185 ;
		RECT	1.045 213.16 1.175 213.21 ;
		RECT	1.34 213.16 1.47 213.21 ;
		RECT	4.47 213.16 4.6 213.21 ;
		RECT	0.9 213.525 14.055 213.705 ;
		RECT	3.02 214.015 3.15 214.065 ;
		RECT	1.57 214.04 1.62 214.17 ;
		RECT	4.87 214.04 4.92 214.17 ;
		RECT	6.375 214.04 6.425 214.17 ;
		RECT	7.015 214.04 7.065 214.17 ;
		RECT	10.27 214.04 10.32 214.17 ;
		RECT	12.79 214.04 12.84 214.17 ;
		RECT	14.33 214.04 14.38 214.17 ;
		RECT	3.02 214.145 3.15 214.195 ;
		RECT	4.035 214.535 4.085 214.665 ;
		RECT	12.655 214.535 12.705 214.665 ;
		RECT	13.9 214.535 13.95 214.665 ;
		RECT	3.02 215 3.15 215.05 ;
		RECT	1.57 215.025 1.62 215.155 ;
		RECT	4.87 215.025 4.92 215.155 ;
		RECT	6.375 215.025 6.425 215.155 ;
		RECT	7.015 215.025 7.065 215.155 ;
		RECT	10.27 215.025 10.32 215.155 ;
		RECT	12.79 215.025 12.84 215.155 ;
		RECT	14.33 215.025 14.38 215.155 ;
		RECT	3.02 215.13 3.15 215.18 ;
		RECT	6.85 215.31 6.9 215.36 ;
		RECT	4.035 215.515 4.085 215.645 ;
		RECT	12.655 215.515 12.705 215.645 ;
		RECT	3.02 215.985 3.15 216.035 ;
		RECT	1.57 216.01 1.62 216.14 ;
		RECT	4.87 216.01 4.92 216.14 ;
		RECT	6.375 216.01 6.425 216.14 ;
		RECT	10.27 216.01 10.32 216.14 ;
		RECT	12.79 216.01 12.84 216.14 ;
		RECT	14.33 216.01 14.38 216.14 ;
		RECT	3.02 216.115 3.15 216.165 ;
		RECT	3.8 216.475 3.93 216.525 ;
		RECT	5.635 216.475 5.765 216.525 ;
		RECT	8.31 216.475 8.44 216.525 ;
		RECT	8.73 216.475 8.86 216.525 ;
		RECT	0.9 216.5 0.95 216.63 ;
		RECT	2.485 216.5 2.535 216.63 ;
		RECT	2.615 216.5 2.665 216.63 ;
		RECT	6.065 216.5 6.115 216.63 ;
		RECT	6.725 216.5 6.775 216.63 ;
		RECT	11.555 216.5 12.57 216.63 ;
		RECT	14.005 216.5 14.055 216.63 ;
		RECT	3.8 216.605 3.93 216.655 ;
		RECT	5.635 216.605 5.765 216.655 ;
		RECT	8.31 216.605 8.44 216.655 ;
		RECT	8.73 216.605 8.86 216.655 ;
		RECT	1.045 216.97 1.175 217.02 ;
		RECT	1.34 216.97 1.47 217.02 ;
		RECT	4.47 216.97 4.6 217.02 ;
		RECT	9.275 216.97 9.405 217.02 ;
		RECT	1.86 216.995 1.91 217.125 ;
		RECT	2.01 216.995 2.06 217.125 ;
		RECT	2.32 216.995 2.37 217.125 ;
		RECT	3.25 216.995 3.3 217.125 ;
		RECT	3.515 216.995 3.565 217.125 ;
		RECT	6.22 216.995 6.27 217.125 ;
		RECT	7.5 216.995 7.55 217.125 ;
		RECT	9.72 216.995 9.77 217.125 ;
		RECT	11.025 216.995 11.075 217.125 ;
		RECT	1.045 217.1 1.175 217.15 ;
		RECT	1.34 217.1 1.47 217.15 ;
		RECT	4.47 217.1 4.6 217.15 ;
		RECT	9.275 217.1 9.405 217.15 ;
		RECT	3.8 217.46 3.93 217.51 ;
		RECT	5.635 217.46 5.765 217.51 ;
		RECT	8.31 217.46 8.44 217.51 ;
		RECT	8.73 217.46 8.86 217.51 ;
		RECT	0.9 217.485 0.95 217.615 ;
		RECT	2.485 217.485 2.535 217.615 ;
		RECT	2.615 217.485 2.665 217.615 ;
		RECT	6.065 217.485 6.115 217.615 ;
		RECT	6.725 217.485 6.775 217.615 ;
		RECT	11.555 217.485 11.865 217.615 ;
		RECT	12.52 217.485 12.57 217.615 ;
		RECT	14.005 217.485 14.055 217.615 ;
		RECT	3.8 217.59 3.93 217.64 ;
		RECT	5.635 217.59 5.765 217.64 ;
		RECT	8.31 217.59 8.44 217.64 ;
		RECT	8.73 217.59 8.86 217.64 ;
		RECT	3.02 217.95 3.15 218 ;
		RECT	1.57 217.975 1.62 218.105 ;
		RECT	4.87 217.975 4.92 218.105 ;
		RECT	6.375 217.975 6.425 218.105 ;
		RECT	10.27 217.975 10.32 218.105 ;
		RECT	12.79 217.975 12.84 218.105 ;
		RECT	14.33 217.975 14.38 218.105 ;
		RECT	3.02 218.08 3.15 218.13 ;
		RECT	0.9 218.445 14.055 218.625 ;
		RECT	3.02 218.935 3.15 218.985 ;
		RECT	1.57 218.96 1.62 219.09 ;
		RECT	4.87 218.96 4.92 219.09 ;
		RECT	6.375 218.96 6.425 219.09 ;
		RECT	10.27 218.96 10.32 219.09 ;
		RECT	12.79 218.96 12.84 219.09 ;
		RECT	14.33 218.96 14.38 219.09 ;
		RECT	3.02 219.065 3.15 219.115 ;
		RECT	12.655 219.445 12.705 219.575 ;
		RECT	4.035 219.455 4.085 219.585 ;
		RECT	3.02 219.92 3.15 219.97 ;
		RECT	1.57 219.945 1.62 220.075 ;
		RECT	4.87 219.945 4.92 220.075 ;
		RECT	6.375 219.945 6.425 220.075 ;
		RECT	10.27 219.945 10.32 220.075 ;
		RECT	12.79 219.945 12.84 220.075 ;
		RECT	14.33 219.945 14.38 220.075 ;
		RECT	3.02 220.05 3.15 220.1 ;
		RECT	0.9 220.41 14.055 220.59 ;
		RECT	14.29 220.72 14.42 220.77 ;
		RECT	1.045 220.905 1.175 220.955 ;
		RECT	1.34 220.905 1.47 220.955 ;
		RECT	4.47 220.905 4.6 220.955 ;
		RECT	9.275 220.905 9.405 220.955 ;
		RECT	1.86 220.93 1.91 221.06 ;
		RECT	2.01 220.93 2.06 221.06 ;
		RECT	2.32 220.93 2.37 221.06 ;
		RECT	3.25 220.93 3.3 221.06 ;
		RECT	3.515 220.93 3.565 221.06 ;
		RECT	6.22 220.93 6.27 221.06 ;
		RECT	7.5 220.93 7.55 221.06 ;
		RECT	9.72 220.93 9.77 221.06 ;
		RECT	11.025 220.93 11.075 221.06 ;
		RECT	1.045 221.035 1.175 221.085 ;
		RECT	1.34 221.035 1.47 221.085 ;
		RECT	4.47 221.035 4.6 221.085 ;
		RECT	9.275 221.035 9.405 221.085 ;
		RECT	0.9 221.215 0.95 221.265 ;
		RECT	2.51 221.215 2.64 221.265 ;
		RECT	0.9 221.395 14.055 221.575 ;
		RECT	2.18 221.915 2.23 222.045 ;
		RECT	8.56 221.915 8.61 222.045 ;
		RECT	10.27 221.915 10.32 222.045 ;
		RECT	4.035 222.405 4.085 222.535 ;
		RECT	3.02 222.87 3.15 222.92 ;
		RECT	1.57 222.895 1.62 223.025 ;
		RECT	4.87 222.895 4.92 223.025 ;
		RECT	6.375 222.895 6.425 223.025 ;
		RECT	11.69 222.895 11.74 223.025 ;
		RECT	12.79 222.895 12.84 223.025 ;
		RECT	12.79 222.895 12.84 223.025 ;
		RECT	14.33 222.895 14.38 223.025 ;
		RECT	3.02 223 3.15 223.05 ;
		RECT	4.035 223.355 4.085 223.485 ;
		RECT	12.655 223.355 12.705 223.485 ;
		RECT	3.02 223.855 3.15 223.905 ;
		RECT	1.57 223.88 1.62 224.01 ;
		RECT	4.87 223.88 4.92 224.01 ;
		RECT	6.375 223.88 6.425 224.01 ;
		RECT	11.69 223.88 11.74 224.01 ;
		RECT	12.79 223.88 12.84 224.01 ;
		RECT	12.79 223.88 12.84 224.01 ;
		RECT	14.33 223.88 14.38 224.01 ;
		RECT	3.02 223.985 3.15 224.035 ;
		RECT	0.9 224.315 14.055 224.495 ;
		RECT	1.045 224.855 1.175 224.905 ;
		RECT	1.34 224.855 1.47 224.905 ;
		RECT	4.47 224.855 4.6 224.905 ;
		RECT	9.275 224.855 9.405 224.905 ;
		RECT	1.86 224.88 1.91 225.01 ;
		RECT	2.01 224.88 2.06 225.01 ;
		RECT	3.25 224.88 3.3 225.01 ;
		RECT	3.515 224.88 3.565 225.01 ;
		RECT	6.22 224.88 6.27 225.01 ;
		RECT	7.5 224.88 7.55 225.01 ;
		RECT	9.72 224.88 9.77 225.01 ;
		RECT	11.025 224.88 11.075 225.01 ;
		RECT	1.045 224.985 1.175 225.035 ;
		RECT	1.34 224.985 1.47 225.035 ;
		RECT	4.47 224.985 4.6 225.035 ;
		RECT	9.275 224.985 9.405 225.035 ;
		RECT	12.655 225.155 12.705 225.205 ;
		RECT	1.045 225.33 1.175 225.38 ;
		RECT	1.34 225.33 1.47 225.38 ;
		RECT	4.47 225.33 4.6 225.38 ;
		RECT	9.275 225.33 9.405 225.38 ;
		RECT	1.86 225.355 1.91 225.485 ;
		RECT	2.01 225.355 2.06 225.485 ;
		RECT	3.25 225.355 3.3 225.485 ;
		RECT	3.515 225.355 3.565 225.485 ;
		RECT	6.22 225.355 6.27 225.485 ;
		RECT	7.5 225.355 7.55 225.485 ;
		RECT	9.72 225.355 9.77 225.485 ;
		RECT	11.025 225.355 11.075 225.485 ;
		RECT	13.675 225.355 13.725 225.485 ;
		RECT	1.045 225.46 1.175 225.51 ;
		RECT	1.34 225.46 1.47 225.51 ;
		RECT	4.47 225.46 4.6 225.51 ;
		RECT	9.275 225.46 9.405 225.51 ;
		RECT	3.02 225.825 3.15 225.875 ;
		RECT	1.57 225.85 1.62 225.98 ;
		RECT	4.87 225.85 4.92 225.98 ;
		RECT	6.375 225.85 6.425 225.98 ;
		RECT	8.975 225.85 9.025 225.98 ;
		RECT	11.69 225.85 11.74 225.98 ;
		RECT	12.79 225.85 12.84 225.98 ;
		RECT	14.33 225.85 14.38 225.98 ;
		RECT	3.02 225.955 3.15 226.005 ;
		RECT	12.655 226.135 12.705 226.185 ;
		RECT	0.9 226.315 14.055 226.495 ;
		RECT	1.57 226.835 1.62 226.965 ;
		RECT	4.87 226.835 4.92 226.965 ;
		RECT	6.375 226.835 6.425 226.965 ;
		RECT	8.975 226.835 9.025 226.965 ;
		RECT	11.69 226.835 11.74 226.965 ;
		RECT	12.79 226.835 12.84 226.965 ;
		RECT	14.33 226.835 14.38 226.965 ;
		RECT	3.02 226.875 3.15 226.925 ;
		RECT	1.045 227.12 1.175 227.17 ;
		RECT	1.34 227.12 1.47 227.17 ;
		RECT	4.47 227.12 4.6 227.17 ;
		RECT	9.275 227.12 9.405 227.17 ;
		RECT	1.86 227.145 1.91 227.275 ;
		RECT	2.01 227.145 2.06 227.275 ;
		RECT	3.25 227.145 3.3 227.275 ;
		RECT	3.515 227.145 3.565 227.275 ;
		RECT	6.22 227.145 6.27 227.275 ;
		RECT	7.5 227.145 7.55 227.275 ;
		RECT	9.72 227.145 9.77 227.275 ;
		RECT	11.025 227.145 11.075 227.275 ;
		RECT	1.045 227.25 1.175 227.3 ;
		RECT	1.34 227.25 1.47 227.3 ;
		RECT	4.47 227.25 4.6 227.3 ;
		RECT	9.275 227.25 9.405 227.3 ;
		RECT	13.8 227.625 13.85 227.755 ;
		RECT	2.18 227.855 2.23 227.985 ;
		RECT	8.56 227.855 8.61 227.985 ;
		RECT	10.27 227.855 10.32 227.985 ;
		RECT	0.62 228.085 0.67 228.215 ;
		RECT	3.65 228.085 3.7 228.215 ;
		RECT	7.19 228.085 7.24 228.215 ;
		RECT	14.14 228.085 14.19 228.215 ;
		RECT	1.085 228.315 1.135 228.445 ;
		RECT	1.38 228.315 1.43 228.445 ;
		RECT	1.86 228.315 1.91 228.445 ;
		RECT	2.01 228.315 2.06 228.445 ;
		RECT	3.25 228.315 3.3 228.445 ;
		RECT	3.515 228.315 3.565 228.445 ;
		RECT	4.51 228.315 4.56 228.445 ;
		RECT	6.22 228.315 6.27 228.445 ;
		RECT	7.5 228.315 7.55 228.445 ;
		RECT	9.315 228.315 9.365 228.445 ;
		RECT	9.72 228.315 9.77 228.445 ;
		RECT	11.025 228.315 11.075 228.445 ;
		RECT	0.435 187.965 0.485 188.095 ;
		RECT	0.435 188.945 0.485 189.075 ;
		RECT	0.435 190.915 0.485 191.045 ;
		RECT	0.435 191.9 0.485 192.03 ;
		RECT	0.435 194.855 0.485 194.985 ;
		RECT	0.435 195.835 0.485 195.965 ;
		RECT	0.435 196.82 0.485 196.95 ;
		RECT	0.435 198.79 0.485 198.92 ;
		RECT	0.17 199.57 0.22 199.62 ;
		RECT	0.435 199.77 0.485 199.9 ;
		RECT	0.435 200.755 0.485 200.885 ;
		RECT	0.18 201.535 0.23 201.585 ;
		RECT	0.435 202.73 0.485 202.86 ;
		RECT	0.435 203.71 0.485 203.84 ;
		RECT	0.435 206.66 0.485 206.79 ;
		RECT	0.435 208.135 0.485 208.265 ;
		RECT	0.435 211.085 0.485 211.215 ;
		RECT	0.435 212.075 0.485 212.205 ;
		RECT	0.18 212.85 0.23 212.9 ;
		RECT	0.435 214.04 0.485 214.17 ;
		RECT	0.435 215.025 0.485 215.155 ;
		RECT	0.17 215.31 0.22 215.36 ;
		RECT	0.435 216.01 0.485 216.14 ;
		RECT	0.435 217.975 0.485 218.105 ;
		RECT	0.435 218.96 0.485 219.09 ;
		RECT	0.435 219.945 0.485 220.075 ;
		RECT	0.17 221.215 0.22 221.265 ;
		RECT	0.435 222.2 0.485 222.25 ;
		RECT	0.435 222.69 0.485 222.74 ;
		RECT	0.435 222.895 0.485 223.025 ;
		RECT	0.435 223.88 0.485 224.01 ;
		RECT	0.435 225.85 0.485 225.98 ;
		RECT	0.435 226.835 0.485 226.965 ;
		RECT	1.57 186.415 1.62 186.545 ;
		RECT	3.06 186.415 3.11 186.545 ;
		RECT	4.87 186.415 4.92 186.545 ;
		RECT	12.79 186.415 12.84 186.545 ;
		RECT	1.57 187.58 1.62 187.71 ;
		RECT	3.02 187.555 3.15 187.735 ;
		RECT	4.87 187.58 4.92 187.71 ;
		RECT	8.955 187.58 9.005 187.71 ;
		RECT	12.79 187.58 12.84 187.71 ;
		RECT	14.29 187.555 14.42 187.735 ;
		RECT	1.045 187.94 1.175 188.12 ;
		RECT	1.34 187.94 1.47 188.12 ;
		RECT	1.86 187.965 1.91 188.095 ;
		RECT	2.01 187.965 2.06 188.095 ;
		RECT	3.25 187.965 3.3 188.095 ;
		RECT	3.515 187.965 3.565 188.095 ;
		RECT	4.47 187.94 4.6 188.12 ;
		RECT	5.035 187.965 5.085 188.095 ;
		RECT	6.22 187.965 6.27 188.095 ;
		RECT	7.5 187.965 7.55 188.095 ;
		RECT	9.275 187.94 9.405 188.12 ;
		RECT	9.72 187.965 9.77 188.095 ;
		RECT	11.025 187.965 11.075 188.095 ;
		RECT	1.045 188.92 1.175 189.1 ;
		RECT	1.34 188.92 1.47 189.1 ;
		RECT	1.86 188.945 1.91 189.075 ;
		RECT	2.01 188.945 2.06 189.075 ;
		RECT	3.25 188.945 3.3 189.075 ;
		RECT	3.515 188.945 3.565 189.075 ;
		RECT	4.47 188.92 4.6 189.1 ;
		RECT	5.035 188.945 5.085 189.075 ;
		RECT	6.22 188.945 6.27 189.075 ;
		RECT	7.5 188.945 7.55 189.075 ;
		RECT	9.275 188.92 9.405 189.1 ;
		RECT	9.72 188.945 9.77 189.075 ;
		RECT	11.025 188.945 11.075 189.075 ;
		RECT	1.57 189.445 1.62 189.575 ;
		RECT	3.02 189.42 3.15 189.6 ;
		RECT	4.87 189.445 4.92 189.575 ;
		RECT	5.9 189.445 5.95 189.575 ;
		RECT	8.955 189.445 9.005 189.575 ;
		RECT	1.57 189.915 1.62 190.045 ;
		RECT	3.02 189.89 3.15 190.07 ;
		RECT	4.87 189.915 4.92 190.045 ;
		RECT	5.9 189.915 5.95 190.045 ;
		RECT	8.955 189.915 9.005 190.045 ;
		RECT	12.79 189.915 12.84 190.045 ;
		RECT	1.045 190.89 1.175 191.07 ;
		RECT	1.34 190.89 1.47 191.07 ;
		RECT	1.86 190.915 1.91 191.045 ;
		RECT	2.01 190.915 2.06 191.045 ;
		RECT	3.25 190.915 3.3 191.045 ;
		RECT	3.515 190.915 3.565 191.045 ;
		RECT	4.47 190.89 4.6 191.07 ;
		RECT	5.035 190.915 5.085 191.045 ;
		RECT	6.22 190.915 6.27 191.045 ;
		RECT	7.5 190.915 7.55 191.045 ;
		RECT	9.275 190.89 9.405 191.07 ;
		RECT	9.72 190.915 9.77 191.045 ;
		RECT	11.025 190.915 11.075 191.045 ;
		RECT	1.045 191.875 1.175 192.055 ;
		RECT	1.34 191.875 1.47 192.055 ;
		RECT	1.86 191.9 1.91 192.03 ;
		RECT	2.01 191.9 2.06 192.03 ;
		RECT	3.25 191.9 3.3 192.03 ;
		RECT	3.515 191.9 3.565 192.03 ;
		RECT	4.47 191.875 4.6 192.055 ;
		RECT	5.035 191.9 5.085 192.03 ;
		RECT	6.22 191.9 6.27 192.03 ;
		RECT	7.5 191.9 7.55 192.03 ;
		RECT	9.72 191.9 9.77 192.03 ;
		RECT	11.025 191.9 11.075 192.03 ;
		RECT	1.57 193.87 1.62 194 ;
		RECT	3.02 193.845 3.15 194.025 ;
		RECT	4.87 193.87 4.92 194 ;
		RECT	5.9 193.87 5.95 194 ;
		RECT	12.79 193.87 12.84 194 ;
		RECT	14.29 193.845 14.42 194.025 ;
		RECT	1.045 194.83 1.175 195.01 ;
		RECT	1.34 194.83 1.47 195.01 ;
		RECT	1.86 194.855 1.91 194.985 ;
		RECT	2.01 194.855 2.06 194.985 ;
		RECT	2.32 194.855 2.37 194.985 ;
		RECT	3.25 194.855 3.3 194.985 ;
		RECT	3.515 194.855 3.565 194.985 ;
		RECT	4.47 194.83 4.6 195.01 ;
		RECT	5.035 194.855 5.085 194.985 ;
		RECT	6.22 194.855 6.27 194.985 ;
		RECT	7.5 194.855 7.55 194.985 ;
		RECT	9.72 194.855 9.77 194.985 ;
		RECT	11.025 194.855 11.075 194.985 ;
		RECT	1.045 195.81 1.175 195.99 ;
		RECT	1.34 195.81 1.47 195.99 ;
		RECT	1.86 195.835 1.91 195.965 ;
		RECT	2.01 195.835 2.06 195.965 ;
		RECT	2.32 195.835 2.37 195.965 ;
		RECT	3.25 195.835 3.3 195.965 ;
		RECT	3.515 195.835 3.565 195.965 ;
		RECT	4.47 195.81 4.6 195.99 ;
		RECT	5.035 195.835 5.085 195.965 ;
		RECT	6.22 195.835 6.27 195.965 ;
		RECT	7.5 195.835 7.55 195.965 ;
		RECT	9.72 195.835 9.77 195.965 ;
		RECT	11.025 195.835 11.075 195.965 ;
		RECT	1.045 196.795 1.175 196.975 ;
		RECT	1.34 196.795 1.47 196.975 ;
		RECT	1.86 196.82 1.91 196.95 ;
		RECT	2.01 196.82 2.06 196.95 ;
		RECT	2.32 196.82 2.37 196.95 ;
		RECT	3.25 196.82 3.3 196.95 ;
		RECT	3.515 196.82 3.565 196.95 ;
		RECT	4.47 196.795 4.6 196.975 ;
		RECT	5.035 196.82 5.085 196.95 ;
		RECT	6.22 196.82 6.27 196.95 ;
		RECT	7.5 196.82 7.55 196.95 ;
		RECT	9.72 196.82 9.77 196.95 ;
		RECT	11.025 196.82 11.075 196.95 ;
		RECT	1.57 197.805 1.62 197.935 ;
		RECT	3.02 197.78 3.15 197.96 ;
		RECT	4.87 197.805 4.92 197.935 ;
		RECT	5.9 197.805 5.95 197.935 ;
		RECT	9.43 197.805 9.48 197.935 ;
		RECT	10.27 197.805 10.32 197.935 ;
		RECT	12.79 197.805 12.84 197.935 ;
		RECT	14.29 197.78 14.42 197.96 ;
		RECT	1.045 198.765 1.175 198.945 ;
		RECT	1.34 198.765 1.47 198.945 ;
		RECT	1.86 198.79 1.91 198.92 ;
		RECT	2.01 198.79 2.06 198.92 ;
		RECT	2.32 198.79 2.37 198.92 ;
		RECT	3.25 198.79 3.3 198.92 ;
		RECT	3.515 198.79 3.565 198.92 ;
		RECT	4.47 198.765 4.6 198.945 ;
		RECT	5.035 198.79 5.085 198.92 ;
		RECT	6.22 198.79 6.27 198.92 ;
		RECT	7.5 198.79 7.55 198.92 ;
		RECT	9.72 198.79 9.77 198.92 ;
		RECT	11.025 198.79 11.075 198.92 ;
		RECT	1.045 199.745 1.175 199.925 ;
		RECT	1.34 199.745 1.47 199.925 ;
		RECT	1.86 199.77 1.91 199.9 ;
		RECT	2.01 199.77 2.06 199.9 ;
		RECT	2.32 199.77 2.37 199.9 ;
		RECT	3.25 199.77 3.3 199.9 ;
		RECT	3.515 199.77 3.565 199.9 ;
		RECT	4.47 199.745 4.6 199.925 ;
		RECT	5.035 199.77 5.085 199.9 ;
		RECT	6.22 199.77 6.27 199.9 ;
		RECT	7.5 199.77 7.55 199.9 ;
		RECT	9.72 199.77 9.77 199.9 ;
		RECT	11.025 199.77 11.075 199.9 ;
		RECT	1.045 200.73 1.175 200.91 ;
		RECT	1.34 200.73 1.47 200.91 ;
		RECT	1.86 200.755 1.91 200.885 ;
		RECT	2.01 200.755 2.06 200.885 ;
		RECT	2.32 200.755 2.37 200.885 ;
		RECT	3.25 200.755 3.3 200.885 ;
		RECT	3.515 200.755 3.565 200.885 ;
		RECT	4.47 200.73 4.6 200.91 ;
		RECT	5.035 200.755 5.085 200.885 ;
		RECT	6.22 200.755 6.27 200.885 ;
		RECT	7.5 200.755 7.55 200.885 ;
		RECT	9.72 200.755 9.77 200.885 ;
		RECT	11.025 200.755 11.075 200.885 ;
		RECT	1.57 201.74 1.62 201.87 ;
		RECT	3.02 201.715 3.15 201.895 ;
		RECT	4.87 201.74 4.92 201.87 ;
		RECT	5.9 201.74 5.95 201.87 ;
		RECT	6.375 201.74 6.425 201.87 ;
		RECT	7.015 201.74 7.065 201.87 ;
		RECT	10.27 201.74 10.32 201.87 ;
		RECT	12.79 201.74 12.84 201.87 ;
		RECT	14.29 201.715 14.42 201.895 ;
		RECT	1.045 202.705 1.175 202.885 ;
		RECT	1.34 202.705 1.47 202.885 ;
		RECT	1.86 202.73 1.91 202.86 ;
		RECT	2.01 202.73 2.06 202.86 ;
		RECT	2.32 202.73 2.37 202.86 ;
		RECT	3.25 202.73 3.3 202.86 ;
		RECT	3.515 202.73 3.565 202.86 ;
		RECT	4.47 202.705 4.6 202.885 ;
		RECT	5.035 202.73 5.085 202.86 ;
		RECT	6.22 202.73 6.27 202.86 ;
		RECT	7.5 202.73 7.55 202.86 ;
		RECT	9.72 202.73 9.77 202.86 ;
		RECT	11.025 202.73 11.075 202.86 ;
		RECT	1.045 203.685 1.175 203.865 ;
		RECT	1.34 203.685 1.47 203.865 ;
		RECT	1.86 203.71 1.91 203.84 ;
		RECT	2.01 203.71 2.06 203.84 ;
		RECT	2.32 203.71 2.37 203.84 ;
		RECT	3.25 203.71 3.3 203.84 ;
		RECT	3.515 203.71 3.565 203.84 ;
		RECT	4.47 203.685 4.6 203.865 ;
		RECT	5.035 203.71 5.085 203.84 ;
		RECT	6.22 203.71 6.27 203.84 ;
		RECT	7.5 203.71 7.55 203.84 ;
		RECT	9.72 203.71 9.77 203.84 ;
		RECT	11.025 203.71 11.075 203.84 ;
		RECT	1.57 204.865 1.62 204.995 ;
		RECT	3.06 204.865 3.11 204.995 ;
		RECT	4.87 204.865 4.92 204.995 ;
		RECT	5.9 204.865 5.95 204.995 ;
		RECT	6.375 204.865 6.425 204.995 ;
		RECT	7.015 204.865 7.065 204.995 ;
		RECT	9.11 204.865 9.16 204.995 ;
		RECT	10.27 204.865 10.32 204.995 ;
		RECT	1.57 205.675 1.62 205.805 ;
		RECT	3.02 205.65 3.15 205.83 ;
		RECT	4.87 205.675 4.92 205.805 ;
		RECT	5.9 205.675 5.95 205.805 ;
		RECT	6.375 205.675 6.425 205.805 ;
		RECT	7.015 205.675 7.065 205.805 ;
		RECT	9.11 205.675 9.16 205.805 ;
		RECT	10.27 205.675 10.32 205.805 ;
		RECT	12.79 205.675 12.84 205.805 ;
		RECT	1.045 206.635 1.175 206.815 ;
		RECT	1.34 206.635 1.47 206.815 ;
		RECT	1.86 206.66 1.91 206.79 ;
		RECT	2.01 206.66 2.06 206.79 ;
		RECT	2.32 206.66 2.37 206.79 ;
		RECT	3.25 206.66 3.3 206.79 ;
		RECT	3.515 206.66 3.565 206.79 ;
		RECT	4.47 206.635 4.6 206.815 ;
		RECT	5.035 206.66 5.085 206.79 ;
		RECT	6.22 206.66 6.27 206.79 ;
		RECT	7.5 206.66 7.55 206.79 ;
		RECT	9.72 206.66 9.77 206.79 ;
		RECT	11.025 206.66 11.075 206.79 ;
		RECT	1.045 208.11 1.175 208.29 ;
		RECT	1.34 208.11 1.47 208.29 ;
		RECT	1.86 208.135 1.91 208.265 ;
		RECT	2.01 208.135 2.06 208.265 ;
		RECT	2.32 208.135 2.37 208.265 ;
		RECT	3.25 208.135 3.3 208.265 ;
		RECT	3.515 208.135 3.565 208.265 ;
		RECT	4.47 208.11 4.6 208.29 ;
		RECT	5.035 208.135 5.085 208.265 ;
		RECT	6.22 208.135 6.27 208.265 ;
		RECT	7.5 208.135 7.55 208.265 ;
		RECT	9.72 208.135 9.77 208.265 ;
		RECT	11.025 208.135 11.075 208.265 ;
		RECT	1.57 209.12 1.62 209.25 ;
		RECT	3.02 209.095 3.15 209.275 ;
		RECT	4.87 209.12 4.92 209.25 ;
		RECT	6.375 209.12 6.425 209.25 ;
		RECT	7.015 209.12 7.065 209.25 ;
		RECT	9.11 209.12 9.16 209.25 ;
		RECT	10.27 209.12 10.32 209.25 ;
		RECT	12.79 209.12 12.84 209.25 ;
		RECT	1.57 209.93 1.62 210.06 ;
		RECT	3.06 209.93 3.11 210.06 ;
		RECT	4.87 209.93 4.92 210.06 ;
		RECT	6.375 209.93 6.425 210.06 ;
		RECT	7.015 209.93 7.065 210.06 ;
		RECT	9.11 209.93 9.16 210.06 ;
		RECT	10.27 209.93 10.32 210.06 ;
		RECT	1.045 211.06 1.175 211.24 ;
		RECT	1.34 211.06 1.47 211.24 ;
		RECT	1.86 211.085 1.91 211.215 ;
		RECT	2.01 211.085 2.06 211.215 ;
		RECT	2.32 211.085 2.37 211.215 ;
		RECT	3.25 211.085 3.3 211.215 ;
		RECT	3.515 211.085 3.565 211.215 ;
		RECT	4.47 211.06 4.6 211.24 ;
		RECT	5.035 211.085 5.085 211.215 ;
		RECT	6.22 211.085 6.27 211.215 ;
		RECT	7.5 211.085 7.55 211.215 ;
		RECT	9.72 211.085 9.77 211.215 ;
		RECT	11.025 211.085 11.075 211.215 ;
		RECT	1.045 212.05 1.175 212.23 ;
		RECT	1.34 212.05 1.47 212.23 ;
		RECT	1.86 212.075 1.91 212.205 ;
		RECT	2.01 212.075 2.06 212.205 ;
		RECT	2.32 212.075 2.37 212.205 ;
		RECT	3.25 212.075 3.3 212.205 ;
		RECT	3.515 212.075 3.565 212.205 ;
		RECT	4.47 212.05 4.6 212.23 ;
		RECT	5.035 212.075 5.085 212.205 ;
		RECT	6.22 212.075 6.27 212.205 ;
		RECT	7.5 212.075 7.55 212.205 ;
		RECT	9.72 212.075 9.77 212.205 ;
		RECT	11.025 212.075 11.075 212.205 ;
		RECT	1.57 213.055 1.62 213.185 ;
		RECT	3.02 213.03 3.15 213.21 ;
		RECT	4.87 213.055 4.92 213.185 ;
		RECT	6.375 213.055 6.425 213.185 ;
		RECT	7.015 213.055 7.065 213.185 ;
		RECT	10.27 213.055 10.32 213.185 ;
		RECT	12.79 213.055 12.84 213.185 ;
		RECT	14.29 213.03 14.42 213.21 ;
		RECT	1.045 214.015 1.175 214.195 ;
		RECT	1.34 214.015 1.47 214.195 ;
		RECT	1.86 214.04 1.91 214.17 ;
		RECT	2.01 214.04 2.06 214.17 ;
		RECT	2.32 214.04 2.37 214.17 ;
		RECT	3.25 214.04 3.3 214.17 ;
		RECT	3.515 214.04 3.565 214.17 ;
		RECT	4.47 214.015 4.6 214.195 ;
		RECT	5.035 214.04 5.085 214.17 ;
		RECT	6.22 214.04 6.27 214.17 ;
		RECT	7.5 214.04 7.55 214.17 ;
		RECT	9.275 214.015 9.405 214.195 ;
		RECT	9.72 214.04 9.77 214.17 ;
		RECT	11.025 214.04 11.075 214.17 ;
		RECT	1.045 215 1.175 215.18 ;
		RECT	1.34 215 1.47 215.18 ;
		RECT	1.86 215.025 1.91 215.155 ;
		RECT	2.01 215.025 2.06 215.155 ;
		RECT	2.32 215.025 2.37 215.155 ;
		RECT	3.25 215.025 3.3 215.155 ;
		RECT	3.515 215.025 3.565 215.155 ;
		RECT	4.47 215 4.6 215.18 ;
		RECT	5.035 215.025 5.085 215.155 ;
		RECT	6.22 215.025 6.27 215.155 ;
		RECT	7.5 215.025 7.55 215.155 ;
		RECT	9.275 215 9.405 215.18 ;
		RECT	9.72 215.025 9.77 215.155 ;
		RECT	11.025 215.025 11.075 215.155 ;
		RECT	1.045 215.985 1.175 216.165 ;
		RECT	1.34 215.985 1.47 216.165 ;
		RECT	1.86 216.01 1.91 216.14 ;
		RECT	2.01 216.01 2.06 216.14 ;
		RECT	2.32 216.01 2.37 216.14 ;
		RECT	3.25 216.01 3.3 216.14 ;
		RECT	3.515 216.01 3.565 216.14 ;
		RECT	4.47 215.985 4.6 216.165 ;
		RECT	6.22 216.01 6.27 216.14 ;
		RECT	7.5 216.01 7.55 216.14 ;
		RECT	9.275 215.985 9.405 216.165 ;
		RECT	9.72 216.01 9.77 216.14 ;
		RECT	11.025 216.01 11.075 216.14 ;
		RECT	1.57 216.995 1.62 217.125 ;
		RECT	3.02 216.97 3.15 217.15 ;
		RECT	4.87 216.995 4.92 217.125 ;
		RECT	6.375 216.995 6.425 217.125 ;
		RECT	10 216.995 10.05 217.125 ;
		RECT	10.27 216.995 10.32 217.125 ;
		RECT	12.79 216.995 12.84 217.125 ;
		RECT	14.29 216.97 14.42 217.15 ;
		RECT	1.045 217.95 1.175 218.13 ;
		RECT	1.34 217.95 1.47 218.13 ;
		RECT	1.86 217.975 1.91 218.105 ;
		RECT	2.01 217.975 2.06 218.105 ;
		RECT	2.32 217.975 2.37 218.105 ;
		RECT	3.25 217.975 3.3 218.105 ;
		RECT	3.515 217.975 3.565 218.105 ;
		RECT	4.47 217.95 4.6 218.13 ;
		RECT	6.22 217.975 6.27 218.105 ;
		RECT	7.5 217.975 7.55 218.105 ;
		RECT	9.275 217.95 9.405 218.13 ;
		RECT	9.72 217.975 9.77 218.105 ;
		RECT	11.025 217.975 11.075 218.105 ;
		RECT	1.045 218.935 1.175 219.115 ;
		RECT	1.34 218.935 1.47 219.115 ;
		RECT	1.86 218.96 1.91 219.09 ;
		RECT	2.01 218.96 2.06 219.09 ;
		RECT	2.32 218.96 2.37 219.09 ;
		RECT	3.25 218.96 3.3 219.09 ;
		RECT	3.515 218.96 3.565 219.09 ;
		RECT	4.47 218.935 4.6 219.115 ;
		RECT	6.22 218.96 6.27 219.09 ;
		RECT	7.5 218.96 7.55 219.09 ;
		RECT	9.275 218.935 9.405 219.115 ;
		RECT	9.72 218.96 9.77 219.09 ;
		RECT	11.025 218.96 11.075 219.09 ;
		RECT	1.045 219.92 1.175 220.1 ;
		RECT	1.34 219.92 1.47 220.1 ;
		RECT	1.86 219.945 1.91 220.075 ;
		RECT	2.01 219.945 2.06 220.075 ;
		RECT	2.32 219.945 2.37 220.075 ;
		RECT	3.25 219.945 3.3 220.075 ;
		RECT	3.515 219.945 3.565 220.075 ;
		RECT	4.47 219.92 4.6 220.1 ;
		RECT	6.22 219.945 6.27 220.075 ;
		RECT	7.5 219.945 7.55 220.075 ;
		RECT	9.275 219.92 9.405 220.1 ;
		RECT	9.72 219.945 9.77 220.075 ;
		RECT	11.025 219.945 11.075 220.075 ;
		RECT	1.57 220.93 1.62 221.06 ;
		RECT	3.02 220.905 3.15 221.085 ;
		RECT	4.87 220.93 4.92 221.06 ;
		RECT	6.375 220.93 6.425 221.06 ;
		RECT	12.79 220.93 12.84 221.06 ;
		RECT	14.29 220.905 14.42 221.085 ;
		RECT	1.045 222.87 1.175 223.05 ;
		RECT	1.34 222.87 1.47 223.05 ;
		RECT	1.86 222.895 1.91 223.025 ;
		RECT	2.01 222.895 2.06 223.025 ;
		RECT	2.32 222.895 2.37 223.025 ;
		RECT	3.25 222.895 3.3 223.025 ;
		RECT	3.515 222.895 3.565 223.025 ;
		RECT	4.47 222.87 4.6 223.05 ;
		RECT	6.22 222.895 6.27 223.025 ;
		RECT	7.5 222.895 7.55 223.025 ;
		RECT	9.275 222.87 9.405 223.05 ;
		RECT	9.72 222.895 9.77 223.025 ;
		RECT	11.025 222.895 11.075 223.025 ;
		RECT	1.045 223.855 1.175 224.035 ;
		RECT	1.34 223.855 1.47 224.035 ;
		RECT	1.86 223.88 1.91 224.01 ;
		RECT	2.01 223.88 2.06 224.01 ;
		RECT	2.32 223.88 2.37 224.01 ;
		RECT	3.25 223.88 3.3 224.01 ;
		RECT	3.515 223.88 3.565 224.01 ;
		RECT	4.47 223.855 4.6 224.035 ;
		RECT	6.22 223.88 6.27 224.01 ;
		RECT	7.5 223.88 7.55 224.01 ;
		RECT	9.275 223.855 9.405 224.035 ;
		RECT	9.72 223.88 9.77 224.01 ;
		RECT	11.025 223.88 11.075 224.01 ;
		RECT	1.57 224.88 1.62 225.01 ;
		RECT	3.02 224.855 3.15 225.035 ;
		RECT	4.87 224.88 4.92 225.01 ;
		RECT	6.375 224.88 6.425 225.01 ;
		RECT	11.69 224.88 11.74 225.01 ;
		RECT	12.79 224.88 12.84 225.01 ;
		RECT	1.57 225.355 1.62 225.485 ;
		RECT	3.02 225.33 3.15 225.51 ;
		RECT	4.87 225.355 4.92 225.485 ;
		RECT	6.375 225.355 6.425 225.485 ;
		RECT	1.045 225.825 1.175 226.005 ;
		RECT	1.34 225.825 1.47 226.005 ;
		RECT	1.86 225.85 1.91 225.98 ;
		RECT	2.01 225.85 2.06 225.98 ;
		RECT	3.25 225.85 3.3 225.98 ;
		RECT	3.515 225.85 3.565 225.98 ;
		RECT	4.47 225.825 4.6 226.005 ;
		RECT	6.22 225.85 6.27 225.98 ;
		RECT	7.5 225.85 7.55 225.98 ;
		RECT	9.275 225.825 9.405 226.005 ;
		RECT	9.72 225.85 9.77 225.98 ;
		RECT	11.025 225.85 11.075 225.98 ;
		RECT	1.86 226.835 1.91 226.965 ;
		RECT	2.01 226.835 2.06 226.965 ;
		RECT	3.25 226.835 3.3 226.965 ;
		RECT	3.515 226.835 3.565 226.965 ;
		RECT	6.22 226.835 6.27 226.965 ;
		RECT	7.5 226.835 7.55 226.965 ;
		RECT	9.72 226.835 9.77 226.965 ;
		RECT	11.025 226.835 11.075 226.965 ;
		RECT	1.57 227.145 1.62 227.275 ;
		RECT	3.02 227.12 3.15 227.3 ;
		RECT	4.87 227.145 4.92 227.275 ;
		RECT	6.375 227.145 6.425 227.275 ;
		RECT	8.975 227.145 9.025 227.275 ;
		RECT	12.79 227.145 12.84 227.275 ;
		RECT	14.29 227.12 14.42 227.3 ;
		RECT	3.06 228.315 3.11 228.445 ;
		RECT	4.87 228.315 4.92 228.445 ;
		RECT	6.375 228.315 6.425 228.445 ;
		RECT	8.975 228.315 9.025 228.445 ;
		RECT	12.79 228.315 12.84 228.445 ;
		RECT	0.9 186.645 0.95 186.775 ;
		RECT	2.485 186.645 2.665 186.775 ;
		RECT	3.84 186.645 3.89 186.775 ;
		RECT	5.675 186.645 5.725 186.775 ;
		RECT	6.065 186.645 6.115 186.775 ;
		RECT	6.725 186.645 6.775 186.775 ;
		RECT	8.35 186.645 8.4 186.775 ;
		RECT	8.77 186.645 8.82 186.775 ;
		RECT	11.555 186.645 11.605 186.775 ;
		RECT	11.815 186.645 11.865 186.775 ;
		RECT	12.52 186.645 12.57 186.775 ;
		RECT	14.005 186.645 14.055 186.775 ;
		RECT	0.62 188.455 0.67 188.585 ;
		RECT	3.65 188.455 3.7 188.585 ;
		RECT	7.18 188.455 7.23 188.585 ;
		RECT	14.14 188.455 14.19 188.585 ;
		RECT	0.62 190.46 0.67 190.59 ;
		RECT	3.65 190.46 3.7 190.59 ;
		RECT	7.18 190.46 7.23 190.59 ;
		RECT	14.14 190.46 14.19 190.59 ;
		RECT	0.62 193.375 0.67 193.505 ;
		RECT	3.65 193.375 3.7 193.505 ;
		RECT	7.18 193.375 7.23 193.505 ;
		RECT	14.14 193.375 14.19 193.505 ;
		RECT	0.62 194.36 0.67 194.49 ;
		RECT	3.65 194.36 3.7 194.49 ;
		RECT	7.18 194.36 7.23 194.49 ;
		RECT	14.14 194.36 14.19 194.49 ;
		RECT	0.62 196.33 0.67 196.46 ;
		RECT	3.65 196.33 3.7 196.46 ;
		RECT	7.18 196.33 7.23 196.46 ;
		RECT	14.14 196.33 14.19 196.46 ;
		RECT	0.62 197.31 0.67 197.44 ;
		RECT	3.65 197.31 3.7 197.44 ;
		RECT	7.18 197.31 7.23 197.44 ;
		RECT	14.14 197.31 14.19 197.44 ;
		RECT	0.62 198.295 0.67 198.425 ;
		RECT	3.65 198.295 3.7 198.425 ;
		RECT	7.18 198.295 7.23 198.425 ;
		RECT	14.14 198.295 14.19 198.425 ;
		RECT	0.62 201.25 0.67 201.38 ;
		RECT	3.65 201.25 3.7 201.38 ;
		RECT	7.18 201.25 7.23 201.38 ;
		RECT	14.14 201.25 14.19 201.38 ;
		RECT	0.9 202.235 0.95 202.365 ;
		RECT	2.485 202.235 2.665 202.365 ;
		RECT	3.8 202.21 3.93 202.39 ;
		RECT	5.635 202.21 5.765 202.39 ;
		RECT	6.065 202.235 6.115 202.365 ;
		RECT	6.675 202.235 6.725 202.365 ;
		RECT	8.31 202.21 8.44 202.39 ;
		RECT	8.73 202.21 8.86 202.39 ;
		RECT	11.555 202.235 11.605 202.365 ;
		RECT	11.815 202.235 11.865 202.365 ;
		RECT	12.52 202.235 12.57 202.365 ;
		RECT	14.005 202.235 14.055 202.365 ;
		RECT	0.62 205.185 0.67 205.315 ;
		RECT	3.65 205.185 3.7 205.315 ;
		RECT	7.18 205.185 7.23 205.315 ;
		RECT	14.14 205.185 14.19 205.315 ;
		RECT	0.62 206.17 0.67 206.3 ;
		RECT	3.65 206.17 3.7 206.3 ;
		RECT	7.18 206.17 7.23 206.3 ;
		RECT	14.14 206.17 14.19 206.3 ;
		RECT	8.31 207.44 8.44 207.49 ;
		RECT	8.73 207.44 8.86 207.49 ;
		RECT	10.12 207.44 10.17 207.49 ;
		RECT	11.555 207.44 11.605 207.49 ;
		RECT	11.815 207.44 11.865 207.49 ;
		RECT	12.52 207.44 12.57 207.49 ;
		RECT	0.62 208.63 0.67 208.76 ;
		RECT	3.65 208.63 3.7 208.76 ;
		RECT	7.18 208.63 7.23 208.76 ;
		RECT	12.655 208.63 12.705 208.76 ;
		RECT	14.14 208.63 14.19 208.76 ;
		RECT	0.62 209.61 0.67 209.74 ;
		RECT	3.65 209.61 3.7 209.74 ;
		RECT	7.18 209.61 7.23 209.74 ;
		RECT	14.14 209.61 14.19 209.74 ;
		RECT	0.9 212.565 0.95 212.695 ;
		RECT	2.51 212.54 2.64 212.72 ;
		RECT	3.8 212.54 3.93 212.72 ;
		RECT	5.635 212.54 5.765 212.72 ;
		RECT	6.065 212.565 6.115 212.695 ;
		RECT	6.675 212.565 6.725 212.695 ;
		RECT	8.31 212.54 8.44 212.72 ;
		RECT	8.73 212.54 8.86 212.72 ;
		RECT	11.555 212.565 11.605 212.695 ;
		RECT	11.815 212.565 11.865 212.695 ;
		RECT	12.52 212.565 12.57 212.695 ;
		RECT	14.005 212.565 14.055 212.695 ;
		RECT	0.62 213.55 0.67 213.68 ;
		RECT	3.65 213.55 3.7 213.68 ;
		RECT	7.18 213.55 7.23 213.68 ;
		RECT	14.14 213.55 14.19 213.68 ;
		RECT	0.62 216.5 0.67 216.63 ;
		RECT	3.65 216.5 3.7 216.63 ;
		RECT	7.18 216.5 7.23 216.63 ;
		RECT	14.14 216.5 14.19 216.63 ;
		RECT	0.62 217.485 0.67 217.615 ;
		RECT	3.65 217.485 3.7 217.615 ;
		RECT	7.18 217.485 7.23 217.615 ;
		RECT	14.14 217.485 14.19 217.615 ;
		RECT	0.62 218.47 0.67 218.6 ;
		RECT	3.65 218.47 3.7 218.6 ;
		RECT	7.18 218.47 7.23 218.6 ;
		RECT	14.14 218.47 14.19 218.6 ;
		RECT	0.62 220.435 0.67 220.565 ;
		RECT	3.65 220.435 3.7 220.565 ;
		RECT	7.18 220.435 7.23 220.565 ;
		RECT	14.14 220.435 14.19 220.565 ;
		RECT	0.62 221.215 0.67 221.265 ;
		RECT	0.62 221.42 0.67 221.55 ;
		RECT	3.65 221.42 3.7 221.55 ;
		RECT	7.18 221.42 7.23 221.55 ;
		RECT	14.14 221.42 14.19 221.55 ;
		RECT	0.62 224.34 0.67 224.47 ;
		RECT	3.65 224.34 3.7 224.47 ;
		RECT	7.18 224.34 7.23 224.47 ;
		RECT	14.14 224.34 14.19 224.47 ;
		RECT	0.62 226.34 0.67 226.47 ;
		RECT	3.65 226.34 3.7 226.47 ;
		RECT	7.18 226.34 7.23 226.47 ;
		RECT	14.14 226.34 14.19 226.47 ;
		RECT	0.9 228.085 0.95 228.215 ;
		RECT	2.485 228.085 2.665 228.215 ;
		RECT	3.84 228.085 3.89 228.215 ;
		RECT	5.675 228.085 5.725 228.215 ;
		RECT	6.065 228.085 6.115 228.215 ;
		RECT	6.725 228.085 6.775 228.215 ;
		RECT	8.35 228.085 8.4 228.215 ;
		RECT	8.77 228.085 8.82 228.215 ;
		RECT	11.555 228.085 11.605 228.215 ;
		RECT	11.815 228.085 11.865 228.215 ;
		RECT	12.52 228.085 12.57 228.215 ;
		RECT	14.005 228.085 14.055 228.215 ;
		RECT	1.57 186.875 1.62 187.005 ;
		RECT	3.06 186.875 3.11 187.005 ;
		RECT	4.87 186.875 4.92 187.005 ;
		RECT	12.79 186.875 12.84 187.005 ;
		RECT	14.33 186.875 14.38 187.005 ;
		RECT	2.18 187.965 2.23 188.095 ;
		RECT	8.56 187.965 8.61 188.095 ;
		RECT	10.27 187.965 10.32 188.095 ;
		RECT	2.18 188.945 2.23 189.075 ;
		RECT	8.56 188.945 8.61 189.075 ;
		RECT	10.27 188.945 10.32 189.075 ;
		RECT	2.18 190.915 2.23 191.045 ;
		RECT	8.56 190.915 8.61 191.045 ;
		RECT	10.27 190.915 10.32 191.045 ;
		RECT	2.18 191.9 2.23 192.03 ;
		RECT	8.56 191.9 8.61 192.03 ;
		RECT	10.27 191.9 10.32 192.03 ;
		RECT	1.57 192.885 1.62 193.015 ;
		RECT	3.02 192.86 3.15 193.04 ;
		RECT	4.87 192.885 4.92 193.015 ;
		RECT	5.9 192.885 5.95 193.015 ;
		RECT	12.79 192.885 12.84 193.015 ;
		RECT	14.29 192.86 14.42 193.04 ;
		RECT	2.18 194.855 2.23 194.985 ;
		RECT	8.56 194.855 8.61 194.985 ;
		RECT	2.18 195.835 2.23 195.965 ;
		RECT	8.56 195.835 8.61 195.965 ;
		RECT	2.18 196.82 2.23 196.95 ;
		RECT	8.56 196.82 8.61 196.95 ;
		RECT	2.18 198.79 2.23 198.92 ;
		RECT	8.56 198.79 8.61 198.92 ;
		RECT	2.18 199.77 2.23 199.9 ;
		RECT	8.56 199.77 8.61 199.9 ;
		RECT	2.18 200.755 2.23 200.885 ;
		RECT	8.56 200.755 8.61 200.885 ;
		RECT	2.18 202.73 2.23 202.86 ;
		RECT	8.56 202.73 8.61 202.86 ;
		RECT	2.18 203.71 2.23 203.84 ;
		RECT	8.56 203.71 8.61 203.84 ;
		RECT	2.18 206.66 2.23 206.79 ;
		RECT	8.56 206.66 8.61 206.79 ;
		RECT	2.18 208.135 2.23 208.265 ;
		RECT	8.56 208.135 8.61 208.265 ;
		RECT	2.18 211.085 2.23 211.215 ;
		RECT	8.56 211.085 8.61 211.215 ;
		RECT	2.18 212.075 2.23 212.205 ;
		RECT	8.56 212.075 8.61 212.205 ;
		RECT	2.18 214.04 2.23 214.17 ;
		RECT	8.56 214.04 8.61 214.17 ;
		RECT	2.18 215.025 2.23 215.155 ;
		RECT	8.56 215.025 8.61 215.155 ;
		RECT	2.18 216.01 2.23 216.14 ;
		RECT	8.56 216.01 8.61 216.14 ;
		RECT	2.18 217.975 2.23 218.105 ;
		RECT	8.56 217.975 8.61 218.105 ;
		RECT	2.18 218.96 2.23 219.09 ;
		RECT	8.56 218.96 8.61 219.09 ;
		RECT	2.18 219.945 2.23 220.075 ;
		RECT	8.56 219.945 8.61 220.075 ;
		RECT	1.57 221.915 1.62 222.045 ;
		RECT	3.02 221.89 3.15 222.07 ;
		RECT	4.87 221.915 4.92 222.045 ;
		RECT	6.375 221.915 6.425 222.045 ;
		RECT	12.79 221.915 12.84 222.045 ;
		RECT	14.29 221.89 14.42 222.07 ;
		RECT	2.18 222.895 2.23 223.025 ;
		RECT	8.56 222.895 8.61 223.025 ;
		RECT	10.27 222.895 10.32 223.025 ;
		RECT	2.18 223.88 2.23 224.01 ;
		RECT	8.56 223.88 8.61 224.01 ;
		RECT	10.27 223.88 10.32 224.01 ;
		RECT	2.18 225.85 2.23 225.98 ;
		RECT	8.56 225.85 8.61 225.98 ;
		RECT	10.27 225.85 10.32 225.98 ;
		RECT	2.18 226.835 2.23 226.965 ;
		RECT	8.56 226.835 8.61 226.965 ;
		RECT	10.27 226.835 10.32 226.965 ;
		RECT	3.06 227.855 3.11 227.985 ;
		RECT	4.87 227.855 4.92 227.985 ;
		RECT	6.375 227.855 6.425 227.985 ;
		RECT	8.975 227.855 9.025 227.985 ;
		RECT	12.79 227.855 12.84 227.985 ;
		RECT	14.33 227.855 14.38 227.985 ;
		RECT	20.875 0.425 21.055 0.555 ;
		RECT	14.965 0.655 15.015 0.785 ;
		RECT	19.485 0.655 19.535 0.785 ;
		RECT	14.765 0.655 14.815 0.785 ;
		RECT	19.685 0.655 19.735 0.785 ;
		RECT	20.7 0.425 20.75 0.555 ;
		RECT	20.875 414.305 21.055 414.435 ;
		RECT	14.965 414.075 15.015 414.205 ;
		RECT	19.485 414.075 19.535 414.205 ;
		RECT	14.765 414.075 14.815 414.205 ;
		RECT	19.685 414.075 19.735 414.205 ;
		RECT	20.7 414.305 20.75 414.435 ;
		RECT	14.565 3.305 14.615 3.435 ;
		RECT	19.885 3.305 19.935 3.435 ;
		RECT	14.765 3.535 14.815 3.665 ;
		RECT	14.765 1.115 14.815 1.245 ;
		RECT	19.685 3.535 19.735 3.665 ;
		RECT	19.685 1.115 19.735 1.245 ;
		RECT	14.965 3.535 15.015 3.665 ;
		RECT	14.965 1.115 15.015 1.245 ;
		RECT	19.485 3.535 19.535 3.665 ;
		RECT	19.485 1.115 19.535 1.245 ;
		RECT	14.565 184.745 14.615 184.875 ;
		RECT	19.885 184.745 19.935 184.875 ;
		RECT	14.765 184.975 14.815 185.105 ;
		RECT	14.765 182.555 14.815 182.685 ;
		RECT	19.685 184.975 19.735 185.105 ;
		RECT	19.685 182.555 19.735 182.685 ;
		RECT	14.965 184.975 15.015 185.105 ;
		RECT	14.965 182.555 15.015 182.685 ;
		RECT	19.485 184.975 19.535 185.105 ;
		RECT	19.485 182.555 19.535 182.685 ;
		RECT	14.565 181.865 14.615 181.995 ;
		RECT	19.885 181.865 19.935 181.995 ;
		RECT	14.765 182.095 14.815 182.225 ;
		RECT	14.765 179.675 14.815 179.805 ;
		RECT	19.685 182.095 19.735 182.225 ;
		RECT	19.685 179.675 19.735 179.805 ;
		RECT	14.965 182.095 15.015 182.225 ;
		RECT	14.965 179.675 15.015 179.805 ;
		RECT	19.485 182.095 19.535 182.225 ;
		RECT	19.485 179.675 19.535 179.805 ;
		RECT	14.565 155.945 14.615 156.075 ;
		RECT	19.885 155.945 19.935 156.075 ;
		RECT	14.765 156.175 14.815 156.305 ;
		RECT	14.765 153.755 14.815 153.885 ;
		RECT	19.685 156.175 19.735 156.305 ;
		RECT	19.685 153.755 19.735 153.885 ;
		RECT	14.965 156.175 15.015 156.305 ;
		RECT	14.965 153.755 15.015 153.885 ;
		RECT	19.485 156.175 19.535 156.305 ;
		RECT	19.485 153.755 19.535 153.885 ;
		RECT	14.565 153.065 14.615 153.195 ;
		RECT	19.885 153.065 19.935 153.195 ;
		RECT	14.765 153.295 14.815 153.425 ;
		RECT	14.765 150.875 14.815 151.005 ;
		RECT	19.685 153.295 19.735 153.425 ;
		RECT	19.685 150.875 19.735 151.005 ;
		RECT	14.965 153.295 15.015 153.425 ;
		RECT	14.965 150.875 15.015 151.005 ;
		RECT	19.485 153.295 19.535 153.425 ;
		RECT	19.485 150.875 19.535 151.005 ;
		RECT	14.565 150.185 14.615 150.315 ;
		RECT	19.885 150.185 19.935 150.315 ;
		RECT	14.765 150.415 14.815 150.545 ;
		RECT	14.765 147.995 14.815 148.125 ;
		RECT	19.685 150.415 19.735 150.545 ;
		RECT	19.685 147.995 19.735 148.125 ;
		RECT	14.965 150.415 15.015 150.545 ;
		RECT	14.965 147.995 15.015 148.125 ;
		RECT	19.485 150.415 19.535 150.545 ;
		RECT	19.485 147.995 19.535 148.125 ;
		RECT	14.565 147.305 14.615 147.435 ;
		RECT	19.885 147.305 19.935 147.435 ;
		RECT	14.765 147.535 14.815 147.665 ;
		RECT	14.765 145.115 14.815 145.245 ;
		RECT	19.685 147.535 19.735 147.665 ;
		RECT	19.685 145.115 19.735 145.245 ;
		RECT	14.965 147.535 15.015 147.665 ;
		RECT	14.965 145.115 15.015 145.245 ;
		RECT	19.485 147.535 19.535 147.665 ;
		RECT	19.485 145.115 19.535 145.245 ;
		RECT	14.565 144.425 14.615 144.555 ;
		RECT	19.885 144.425 19.935 144.555 ;
		RECT	14.765 144.655 14.815 144.785 ;
		RECT	14.765 142.235 14.815 142.365 ;
		RECT	19.685 144.655 19.735 144.785 ;
		RECT	19.685 142.235 19.735 142.365 ;
		RECT	14.965 144.655 15.015 144.785 ;
		RECT	14.965 142.235 15.015 142.365 ;
		RECT	19.485 144.655 19.535 144.785 ;
		RECT	19.485 142.235 19.535 142.365 ;
		RECT	14.565 141.545 14.615 141.675 ;
		RECT	19.885 141.545 19.935 141.675 ;
		RECT	14.765 141.775 14.815 141.905 ;
		RECT	14.765 139.355 14.815 139.485 ;
		RECT	19.685 141.775 19.735 141.905 ;
		RECT	19.685 139.355 19.735 139.485 ;
		RECT	14.965 141.775 15.015 141.905 ;
		RECT	14.965 139.355 15.015 139.485 ;
		RECT	19.485 141.775 19.535 141.905 ;
		RECT	19.485 139.355 19.535 139.485 ;
		RECT	14.565 138.665 14.615 138.795 ;
		RECT	19.885 138.665 19.935 138.795 ;
		RECT	14.765 138.895 14.815 139.025 ;
		RECT	14.765 136.475 14.815 136.605 ;
		RECT	19.685 138.895 19.735 139.025 ;
		RECT	19.685 136.475 19.735 136.605 ;
		RECT	14.965 138.895 15.015 139.025 ;
		RECT	14.965 136.475 15.015 136.605 ;
		RECT	19.485 138.895 19.535 139.025 ;
		RECT	19.485 136.475 19.535 136.605 ;
		RECT	14.565 135.785 14.615 135.915 ;
		RECT	19.885 135.785 19.935 135.915 ;
		RECT	14.765 136.015 14.815 136.145 ;
		RECT	14.765 133.595 14.815 133.725 ;
		RECT	19.685 136.015 19.735 136.145 ;
		RECT	19.685 133.595 19.735 133.725 ;
		RECT	14.965 136.015 15.015 136.145 ;
		RECT	14.965 133.595 15.015 133.725 ;
		RECT	19.485 136.015 19.535 136.145 ;
		RECT	19.485 133.595 19.535 133.725 ;
		RECT	14.565 132.905 14.615 133.035 ;
		RECT	19.885 132.905 19.935 133.035 ;
		RECT	14.765 133.135 14.815 133.265 ;
		RECT	14.765 130.715 14.815 130.845 ;
		RECT	19.685 133.135 19.735 133.265 ;
		RECT	19.685 130.715 19.735 130.845 ;
		RECT	14.965 133.135 15.015 133.265 ;
		RECT	14.965 130.715 15.015 130.845 ;
		RECT	19.485 133.135 19.535 133.265 ;
		RECT	19.485 130.715 19.535 130.845 ;
		RECT	14.565 130.025 14.615 130.155 ;
		RECT	19.885 130.025 19.935 130.155 ;
		RECT	14.765 130.255 14.815 130.385 ;
		RECT	14.765 127.835 14.815 127.965 ;
		RECT	19.685 130.255 19.735 130.385 ;
		RECT	19.685 127.835 19.735 127.965 ;
		RECT	14.965 130.255 15.015 130.385 ;
		RECT	14.965 127.835 15.015 127.965 ;
		RECT	19.485 130.255 19.535 130.385 ;
		RECT	19.485 127.835 19.535 127.965 ;
		RECT	14.565 178.985 14.615 179.115 ;
		RECT	19.885 178.985 19.935 179.115 ;
		RECT	14.765 179.215 14.815 179.345 ;
		RECT	14.765 176.795 14.815 176.925 ;
		RECT	19.685 179.215 19.735 179.345 ;
		RECT	19.685 176.795 19.735 176.925 ;
		RECT	14.965 179.215 15.015 179.345 ;
		RECT	14.965 176.795 15.015 176.925 ;
		RECT	19.485 179.215 19.535 179.345 ;
		RECT	19.485 176.795 19.535 176.925 ;
		RECT	14.565 127.145 14.615 127.275 ;
		RECT	19.885 127.145 19.935 127.275 ;
		RECT	14.765 127.375 14.815 127.505 ;
		RECT	14.765 124.955 14.815 125.085 ;
		RECT	19.685 127.375 19.735 127.505 ;
		RECT	19.685 124.955 19.735 125.085 ;
		RECT	14.965 127.375 15.015 127.505 ;
		RECT	14.965 124.955 15.015 125.085 ;
		RECT	19.485 127.375 19.535 127.505 ;
		RECT	19.485 124.955 19.535 125.085 ;
		RECT	14.565 124.265 14.615 124.395 ;
		RECT	19.885 124.265 19.935 124.395 ;
		RECT	14.765 124.495 14.815 124.625 ;
		RECT	14.765 122.075 14.815 122.205 ;
		RECT	19.685 124.495 19.735 124.625 ;
		RECT	19.685 122.075 19.735 122.205 ;
		RECT	14.965 124.495 15.015 124.625 ;
		RECT	14.965 122.075 15.015 122.205 ;
		RECT	19.485 124.495 19.535 124.625 ;
		RECT	19.485 122.075 19.535 122.205 ;
		RECT	14.565 121.385 14.615 121.515 ;
		RECT	19.885 121.385 19.935 121.515 ;
		RECT	14.765 121.615 14.815 121.745 ;
		RECT	14.765 119.195 14.815 119.325 ;
		RECT	19.685 121.615 19.735 121.745 ;
		RECT	19.685 119.195 19.735 119.325 ;
		RECT	14.965 121.615 15.015 121.745 ;
		RECT	14.965 119.195 15.015 119.325 ;
		RECT	19.485 121.615 19.535 121.745 ;
		RECT	19.485 119.195 19.535 119.325 ;
		RECT	14.565 118.505 14.615 118.635 ;
		RECT	19.885 118.505 19.935 118.635 ;
		RECT	14.765 118.735 14.815 118.865 ;
		RECT	14.765 116.315 14.815 116.445 ;
		RECT	19.685 118.735 19.735 118.865 ;
		RECT	19.685 116.315 19.735 116.445 ;
		RECT	14.965 118.735 15.015 118.865 ;
		RECT	14.965 116.315 15.015 116.445 ;
		RECT	19.485 118.735 19.535 118.865 ;
		RECT	19.485 116.315 19.535 116.445 ;
		RECT	14.565 115.625 14.615 115.755 ;
		RECT	19.885 115.625 19.935 115.755 ;
		RECT	14.765 115.855 14.815 115.985 ;
		RECT	14.765 113.435 14.815 113.565 ;
		RECT	19.685 115.855 19.735 115.985 ;
		RECT	19.685 113.435 19.735 113.565 ;
		RECT	14.965 115.855 15.015 115.985 ;
		RECT	14.965 113.435 15.015 113.565 ;
		RECT	19.485 115.855 19.535 115.985 ;
		RECT	19.485 113.435 19.535 113.565 ;
		RECT	14.565 112.745 14.615 112.875 ;
		RECT	19.885 112.745 19.935 112.875 ;
		RECT	14.765 112.975 14.815 113.105 ;
		RECT	14.765 110.555 14.815 110.685 ;
		RECT	19.685 112.975 19.735 113.105 ;
		RECT	19.685 110.555 19.735 110.685 ;
		RECT	14.965 112.975 15.015 113.105 ;
		RECT	14.965 110.555 15.015 110.685 ;
		RECT	19.485 112.975 19.535 113.105 ;
		RECT	19.485 110.555 19.535 110.685 ;
		RECT	14.565 109.865 14.615 109.995 ;
		RECT	19.885 109.865 19.935 109.995 ;
		RECT	14.765 110.095 14.815 110.225 ;
		RECT	14.765 107.675 14.815 107.805 ;
		RECT	19.685 110.095 19.735 110.225 ;
		RECT	19.685 107.675 19.735 107.805 ;
		RECT	14.965 110.095 15.015 110.225 ;
		RECT	14.965 107.675 15.015 107.805 ;
		RECT	19.485 110.095 19.535 110.225 ;
		RECT	19.485 107.675 19.535 107.805 ;
		RECT	14.565 106.985 14.615 107.115 ;
		RECT	19.885 106.985 19.935 107.115 ;
		RECT	14.765 107.215 14.815 107.345 ;
		RECT	14.765 104.795 14.815 104.925 ;
		RECT	19.685 107.215 19.735 107.345 ;
		RECT	19.685 104.795 19.735 104.925 ;
		RECT	14.965 107.215 15.015 107.345 ;
		RECT	14.965 104.795 15.015 104.925 ;
		RECT	19.485 107.215 19.535 107.345 ;
		RECT	19.485 104.795 19.535 104.925 ;
		RECT	14.565 104.105 14.615 104.235 ;
		RECT	19.885 104.105 19.935 104.235 ;
		RECT	14.765 104.335 14.815 104.465 ;
		RECT	14.765 101.915 14.815 102.045 ;
		RECT	19.685 104.335 19.735 104.465 ;
		RECT	19.685 101.915 19.735 102.045 ;
		RECT	14.965 104.335 15.015 104.465 ;
		RECT	14.965 101.915 15.015 102.045 ;
		RECT	19.485 104.335 19.535 104.465 ;
		RECT	19.485 101.915 19.535 102.045 ;
		RECT	14.565 101.225 14.615 101.355 ;
		RECT	19.885 101.225 19.935 101.355 ;
		RECT	14.765 101.455 14.815 101.585 ;
		RECT	14.765 99.035 14.815 99.165 ;
		RECT	19.685 101.455 19.735 101.585 ;
		RECT	19.685 99.035 19.735 99.165 ;
		RECT	14.965 101.455 15.015 101.585 ;
		RECT	14.965 99.035 15.015 99.165 ;
		RECT	19.485 101.455 19.535 101.585 ;
		RECT	19.485 99.035 19.535 99.165 ;
		RECT	14.565 176.105 14.615 176.235 ;
		RECT	19.885 176.105 19.935 176.235 ;
		RECT	14.765 176.335 14.815 176.465 ;
		RECT	14.765 173.915 14.815 174.045 ;
		RECT	19.685 176.335 19.735 176.465 ;
		RECT	19.685 173.915 19.735 174.045 ;
		RECT	14.965 176.335 15.015 176.465 ;
		RECT	14.965 173.915 15.015 174.045 ;
		RECT	19.485 176.335 19.535 176.465 ;
		RECT	19.485 173.915 19.535 174.045 ;
		RECT	14.565 98.345 14.615 98.475 ;
		RECT	19.885 98.345 19.935 98.475 ;
		RECT	14.765 98.575 14.815 98.705 ;
		RECT	14.765 96.155 14.815 96.285 ;
		RECT	19.685 98.575 19.735 98.705 ;
		RECT	19.685 96.155 19.735 96.285 ;
		RECT	14.965 98.575 15.015 98.705 ;
		RECT	14.965 96.155 15.015 96.285 ;
		RECT	19.485 98.575 19.535 98.705 ;
		RECT	19.485 96.155 19.535 96.285 ;
		RECT	14.565 95.465 14.615 95.595 ;
		RECT	19.885 95.465 19.935 95.595 ;
		RECT	14.765 95.695 14.815 95.825 ;
		RECT	14.765 93.275 14.815 93.405 ;
		RECT	19.685 95.695 19.735 95.825 ;
		RECT	19.685 93.275 19.735 93.405 ;
		RECT	14.965 95.695 15.015 95.825 ;
		RECT	14.965 93.275 15.015 93.405 ;
		RECT	19.485 95.695 19.535 95.825 ;
		RECT	19.485 93.275 19.535 93.405 ;
		RECT	14.565 92.585 14.615 92.715 ;
		RECT	19.885 92.585 19.935 92.715 ;
		RECT	14.765 92.815 14.815 92.945 ;
		RECT	14.765 90.395 14.815 90.525 ;
		RECT	19.685 92.815 19.735 92.945 ;
		RECT	19.685 90.395 19.735 90.525 ;
		RECT	14.965 92.815 15.015 92.945 ;
		RECT	14.965 90.395 15.015 90.525 ;
		RECT	19.485 92.815 19.535 92.945 ;
		RECT	19.485 90.395 19.535 90.525 ;
		RECT	14.565 89.705 14.615 89.835 ;
		RECT	19.885 89.705 19.935 89.835 ;
		RECT	14.765 89.935 14.815 90.065 ;
		RECT	14.765 87.515 14.815 87.645 ;
		RECT	19.685 89.935 19.735 90.065 ;
		RECT	19.685 87.515 19.735 87.645 ;
		RECT	14.965 89.935 15.015 90.065 ;
		RECT	14.965 87.515 15.015 87.645 ;
		RECT	19.485 89.935 19.535 90.065 ;
		RECT	19.485 87.515 19.535 87.645 ;
		RECT	14.565 86.825 14.615 86.955 ;
		RECT	19.885 86.825 19.935 86.955 ;
		RECT	14.765 87.055 14.815 87.185 ;
		RECT	14.765 84.635 14.815 84.765 ;
		RECT	19.685 87.055 19.735 87.185 ;
		RECT	19.685 84.635 19.735 84.765 ;
		RECT	14.965 87.055 15.015 87.185 ;
		RECT	14.965 84.635 15.015 84.765 ;
		RECT	19.485 87.055 19.535 87.185 ;
		RECT	19.485 84.635 19.535 84.765 ;
		RECT	14.565 83.945 14.615 84.075 ;
		RECT	19.885 83.945 19.935 84.075 ;
		RECT	14.765 84.175 14.815 84.305 ;
		RECT	14.765 81.755 14.815 81.885 ;
		RECT	19.685 84.175 19.735 84.305 ;
		RECT	19.685 81.755 19.735 81.885 ;
		RECT	14.965 84.175 15.015 84.305 ;
		RECT	14.965 81.755 15.015 81.885 ;
		RECT	19.485 84.175 19.535 84.305 ;
		RECT	19.485 81.755 19.535 81.885 ;
		RECT	14.565 81.065 14.615 81.195 ;
		RECT	19.885 81.065 19.935 81.195 ;
		RECT	14.765 81.295 14.815 81.425 ;
		RECT	14.765 78.875 14.815 79.005 ;
		RECT	19.685 81.295 19.735 81.425 ;
		RECT	19.685 78.875 19.735 79.005 ;
		RECT	14.965 81.295 15.015 81.425 ;
		RECT	14.965 78.875 15.015 79.005 ;
		RECT	19.485 81.295 19.535 81.425 ;
		RECT	19.485 78.875 19.535 79.005 ;
		RECT	14.565 78.185 14.615 78.315 ;
		RECT	19.885 78.185 19.935 78.315 ;
		RECT	14.765 78.415 14.815 78.545 ;
		RECT	14.765 75.995 14.815 76.125 ;
		RECT	19.685 78.415 19.735 78.545 ;
		RECT	19.685 75.995 19.735 76.125 ;
		RECT	14.965 78.415 15.015 78.545 ;
		RECT	14.965 75.995 15.015 76.125 ;
		RECT	19.485 78.415 19.535 78.545 ;
		RECT	19.485 75.995 19.535 76.125 ;
		RECT	14.565 75.305 14.615 75.435 ;
		RECT	19.885 75.305 19.935 75.435 ;
		RECT	14.765 75.535 14.815 75.665 ;
		RECT	14.765 73.115 14.815 73.245 ;
		RECT	19.685 75.535 19.735 75.665 ;
		RECT	19.685 73.115 19.735 73.245 ;
		RECT	14.965 75.535 15.015 75.665 ;
		RECT	14.965 73.115 15.015 73.245 ;
		RECT	19.485 75.535 19.535 75.665 ;
		RECT	19.485 73.115 19.535 73.245 ;
		RECT	14.565 72.425 14.615 72.555 ;
		RECT	19.885 72.425 19.935 72.555 ;
		RECT	14.765 72.655 14.815 72.785 ;
		RECT	14.765 70.235 14.815 70.365 ;
		RECT	19.685 72.655 19.735 72.785 ;
		RECT	19.685 70.235 19.735 70.365 ;
		RECT	14.965 72.655 15.015 72.785 ;
		RECT	14.965 70.235 15.015 70.365 ;
		RECT	19.485 72.655 19.535 72.785 ;
		RECT	19.485 70.235 19.535 70.365 ;
		RECT	14.565 173.225 14.615 173.355 ;
		RECT	19.885 173.225 19.935 173.355 ;
		RECT	14.765 173.455 14.815 173.585 ;
		RECT	14.765 171.035 14.815 171.165 ;
		RECT	19.685 173.455 19.735 173.585 ;
		RECT	19.685 171.035 19.735 171.165 ;
		RECT	14.965 173.455 15.015 173.585 ;
		RECT	14.965 171.035 15.015 171.165 ;
		RECT	19.485 173.455 19.535 173.585 ;
		RECT	19.485 171.035 19.535 171.165 ;
		RECT	14.565 69.545 14.615 69.675 ;
		RECT	19.885 69.545 19.935 69.675 ;
		RECT	14.765 69.775 14.815 69.905 ;
		RECT	14.765 67.355 14.815 67.485 ;
		RECT	19.685 69.775 19.735 69.905 ;
		RECT	19.685 67.355 19.735 67.485 ;
		RECT	14.965 69.775 15.015 69.905 ;
		RECT	14.965 67.355 15.015 67.485 ;
		RECT	19.485 69.775 19.535 69.905 ;
		RECT	19.485 67.355 19.535 67.485 ;
		RECT	14.565 66.665 14.615 66.795 ;
		RECT	19.885 66.665 19.935 66.795 ;
		RECT	14.765 66.895 14.815 67.025 ;
		RECT	14.765 64.475 14.815 64.605 ;
		RECT	19.685 66.895 19.735 67.025 ;
		RECT	19.685 64.475 19.735 64.605 ;
		RECT	14.965 66.895 15.015 67.025 ;
		RECT	14.965 64.475 15.015 64.605 ;
		RECT	19.485 66.895 19.535 67.025 ;
		RECT	19.485 64.475 19.535 64.605 ;
		RECT	14.565 63.785 14.615 63.915 ;
		RECT	19.885 63.785 19.935 63.915 ;
		RECT	14.765 64.015 14.815 64.145 ;
		RECT	14.765 61.595 14.815 61.725 ;
		RECT	19.685 64.015 19.735 64.145 ;
		RECT	19.685 61.595 19.735 61.725 ;
		RECT	14.965 64.015 15.015 64.145 ;
		RECT	14.965 61.595 15.015 61.725 ;
		RECT	19.485 64.015 19.535 64.145 ;
		RECT	19.485 61.595 19.535 61.725 ;
		RECT	14.565 60.905 14.615 61.035 ;
		RECT	19.885 60.905 19.935 61.035 ;
		RECT	14.765 61.135 14.815 61.265 ;
		RECT	14.765 58.715 14.815 58.845 ;
		RECT	19.685 61.135 19.735 61.265 ;
		RECT	19.685 58.715 19.735 58.845 ;
		RECT	14.965 61.135 15.015 61.265 ;
		RECT	14.965 58.715 15.015 58.845 ;
		RECT	19.485 61.135 19.535 61.265 ;
		RECT	19.485 58.715 19.535 58.845 ;
		RECT	14.565 58.025 14.615 58.155 ;
		RECT	19.885 58.025 19.935 58.155 ;
		RECT	14.765 58.255 14.815 58.385 ;
		RECT	14.765 55.835 14.815 55.965 ;
		RECT	19.685 58.255 19.735 58.385 ;
		RECT	19.685 55.835 19.735 55.965 ;
		RECT	14.965 58.255 15.015 58.385 ;
		RECT	14.965 55.835 15.015 55.965 ;
		RECT	19.485 58.255 19.535 58.385 ;
		RECT	19.485 55.835 19.535 55.965 ;
		RECT	14.565 55.145 14.615 55.275 ;
		RECT	19.885 55.145 19.935 55.275 ;
		RECT	14.765 55.375 14.815 55.505 ;
		RECT	14.765 52.955 14.815 53.085 ;
		RECT	19.685 55.375 19.735 55.505 ;
		RECT	19.685 52.955 19.735 53.085 ;
		RECT	14.965 55.375 15.015 55.505 ;
		RECT	14.965 52.955 15.015 53.085 ;
		RECT	19.485 55.375 19.535 55.505 ;
		RECT	19.485 52.955 19.535 53.085 ;
		RECT	14.565 52.265 14.615 52.395 ;
		RECT	19.885 52.265 19.935 52.395 ;
		RECT	14.765 52.495 14.815 52.625 ;
		RECT	14.765 50.075 14.815 50.205 ;
		RECT	19.685 52.495 19.735 52.625 ;
		RECT	19.685 50.075 19.735 50.205 ;
		RECT	14.965 52.495 15.015 52.625 ;
		RECT	14.965 50.075 15.015 50.205 ;
		RECT	19.485 52.495 19.535 52.625 ;
		RECT	19.485 50.075 19.535 50.205 ;
		RECT	14.565 49.385 14.615 49.515 ;
		RECT	19.885 49.385 19.935 49.515 ;
		RECT	14.765 49.615 14.815 49.745 ;
		RECT	14.765 47.195 14.815 47.325 ;
		RECT	19.685 49.615 19.735 49.745 ;
		RECT	19.685 47.195 19.735 47.325 ;
		RECT	14.965 49.615 15.015 49.745 ;
		RECT	14.965 47.195 15.015 47.325 ;
		RECT	19.485 49.615 19.535 49.745 ;
		RECT	19.485 47.195 19.535 47.325 ;
		RECT	14.565 46.505 14.615 46.635 ;
		RECT	19.885 46.505 19.935 46.635 ;
		RECT	14.765 46.735 14.815 46.865 ;
		RECT	14.765 44.315 14.815 44.445 ;
		RECT	19.685 46.735 19.735 46.865 ;
		RECT	19.685 44.315 19.735 44.445 ;
		RECT	14.965 46.735 15.015 46.865 ;
		RECT	14.965 44.315 15.015 44.445 ;
		RECT	19.485 46.735 19.535 46.865 ;
		RECT	19.485 44.315 19.535 44.445 ;
		RECT	14.565 43.625 14.615 43.755 ;
		RECT	19.885 43.625 19.935 43.755 ;
		RECT	14.765 43.855 14.815 43.985 ;
		RECT	14.765 41.435 14.815 41.565 ;
		RECT	19.685 43.855 19.735 43.985 ;
		RECT	19.685 41.435 19.735 41.565 ;
		RECT	14.965 43.855 15.015 43.985 ;
		RECT	14.965 41.435 15.015 41.565 ;
		RECT	19.485 43.855 19.535 43.985 ;
		RECT	19.485 41.435 19.535 41.565 ;
		RECT	14.565 170.345 14.615 170.475 ;
		RECT	19.885 170.345 19.935 170.475 ;
		RECT	14.765 170.575 14.815 170.705 ;
		RECT	14.765 168.155 14.815 168.285 ;
		RECT	19.685 170.575 19.735 170.705 ;
		RECT	19.685 168.155 19.735 168.285 ;
		RECT	14.965 170.575 15.015 170.705 ;
		RECT	14.965 168.155 15.015 168.285 ;
		RECT	19.485 170.575 19.535 170.705 ;
		RECT	19.485 168.155 19.535 168.285 ;
		RECT	14.565 40.745 14.615 40.875 ;
		RECT	19.885 40.745 19.935 40.875 ;
		RECT	14.765 40.975 14.815 41.105 ;
		RECT	14.765 38.555 14.815 38.685 ;
		RECT	19.685 40.975 19.735 41.105 ;
		RECT	19.685 38.555 19.735 38.685 ;
		RECT	14.965 40.975 15.015 41.105 ;
		RECT	14.965 38.555 15.015 38.685 ;
		RECT	19.485 40.975 19.535 41.105 ;
		RECT	19.485 38.555 19.535 38.685 ;
		RECT	14.565 37.865 14.615 37.995 ;
		RECT	19.885 37.865 19.935 37.995 ;
		RECT	14.765 38.095 14.815 38.225 ;
		RECT	14.765 35.675 14.815 35.805 ;
		RECT	19.685 38.095 19.735 38.225 ;
		RECT	19.685 35.675 19.735 35.805 ;
		RECT	14.965 38.095 15.015 38.225 ;
		RECT	14.965 35.675 15.015 35.805 ;
		RECT	19.485 38.095 19.535 38.225 ;
		RECT	19.485 35.675 19.535 35.805 ;
		RECT	14.565 34.985 14.615 35.115 ;
		RECT	19.885 34.985 19.935 35.115 ;
		RECT	14.765 35.215 14.815 35.345 ;
		RECT	14.765 32.795 14.815 32.925 ;
		RECT	19.685 35.215 19.735 35.345 ;
		RECT	19.685 32.795 19.735 32.925 ;
		RECT	14.965 35.215 15.015 35.345 ;
		RECT	14.965 32.795 15.015 32.925 ;
		RECT	19.485 35.215 19.535 35.345 ;
		RECT	19.485 32.795 19.535 32.925 ;
		RECT	14.565 32.105 14.615 32.235 ;
		RECT	19.885 32.105 19.935 32.235 ;
		RECT	14.765 32.335 14.815 32.465 ;
		RECT	14.765 29.915 14.815 30.045 ;
		RECT	19.685 32.335 19.735 32.465 ;
		RECT	19.685 29.915 19.735 30.045 ;
		RECT	14.965 32.335 15.015 32.465 ;
		RECT	14.965 29.915 15.015 30.045 ;
		RECT	19.485 32.335 19.535 32.465 ;
		RECT	19.485 29.915 19.535 30.045 ;
		RECT	14.565 29.225 14.615 29.355 ;
		RECT	19.885 29.225 19.935 29.355 ;
		RECT	14.765 29.455 14.815 29.585 ;
		RECT	14.765 27.035 14.815 27.165 ;
		RECT	19.685 29.455 19.735 29.585 ;
		RECT	19.685 27.035 19.735 27.165 ;
		RECT	14.965 29.455 15.015 29.585 ;
		RECT	14.965 27.035 15.015 27.165 ;
		RECT	19.485 29.455 19.535 29.585 ;
		RECT	19.485 27.035 19.535 27.165 ;
		RECT	14.565 26.345 14.615 26.475 ;
		RECT	19.885 26.345 19.935 26.475 ;
		RECT	14.765 26.575 14.815 26.705 ;
		RECT	14.765 24.155 14.815 24.285 ;
		RECT	19.685 26.575 19.735 26.705 ;
		RECT	19.685 24.155 19.735 24.285 ;
		RECT	14.965 26.575 15.015 26.705 ;
		RECT	14.965 24.155 15.015 24.285 ;
		RECT	19.485 26.575 19.535 26.705 ;
		RECT	19.485 24.155 19.535 24.285 ;
		RECT	14.565 23.465 14.615 23.595 ;
		RECT	19.885 23.465 19.935 23.595 ;
		RECT	14.765 23.695 14.815 23.825 ;
		RECT	14.765 21.275 14.815 21.405 ;
		RECT	19.685 23.695 19.735 23.825 ;
		RECT	19.685 21.275 19.735 21.405 ;
		RECT	14.965 23.695 15.015 23.825 ;
		RECT	14.965 21.275 15.015 21.405 ;
		RECT	19.485 23.695 19.535 23.825 ;
		RECT	19.485 21.275 19.535 21.405 ;
		RECT	14.565 20.585 14.615 20.715 ;
		RECT	19.885 20.585 19.935 20.715 ;
		RECT	14.765 20.815 14.815 20.945 ;
		RECT	14.765 18.395 14.815 18.525 ;
		RECT	19.685 20.815 19.735 20.945 ;
		RECT	19.685 18.395 19.735 18.525 ;
		RECT	14.965 20.815 15.015 20.945 ;
		RECT	14.965 18.395 15.015 18.525 ;
		RECT	19.485 20.815 19.535 20.945 ;
		RECT	19.485 18.395 19.535 18.525 ;
		RECT	14.565 17.705 14.615 17.835 ;
		RECT	19.885 17.705 19.935 17.835 ;
		RECT	14.765 17.935 14.815 18.065 ;
		RECT	14.765 15.515 14.815 15.645 ;
		RECT	19.685 17.935 19.735 18.065 ;
		RECT	19.685 15.515 19.735 15.645 ;
		RECT	14.965 17.935 15.015 18.065 ;
		RECT	14.965 15.515 15.015 15.645 ;
		RECT	19.485 17.935 19.535 18.065 ;
		RECT	19.485 15.515 19.535 15.645 ;
		RECT	14.565 14.825 14.615 14.955 ;
		RECT	19.885 14.825 19.935 14.955 ;
		RECT	14.765 15.055 14.815 15.185 ;
		RECT	14.765 12.635 14.815 12.765 ;
		RECT	19.685 15.055 19.735 15.185 ;
		RECT	19.685 12.635 19.735 12.765 ;
		RECT	14.965 15.055 15.015 15.185 ;
		RECT	14.965 12.635 15.015 12.765 ;
		RECT	19.485 15.055 19.535 15.185 ;
		RECT	19.485 12.635 19.535 12.765 ;
		RECT	14.565 167.465 14.615 167.595 ;
		RECT	19.885 167.465 19.935 167.595 ;
		RECT	14.765 167.695 14.815 167.825 ;
		RECT	14.765 165.275 14.815 165.405 ;
		RECT	19.685 167.695 19.735 167.825 ;
		RECT	19.685 165.275 19.735 165.405 ;
		RECT	14.965 167.695 15.015 167.825 ;
		RECT	14.965 165.275 15.015 165.405 ;
		RECT	19.485 167.695 19.535 167.825 ;
		RECT	19.485 165.275 19.535 165.405 ;
		RECT	14.565 11.945 14.615 12.075 ;
		RECT	19.885 11.945 19.935 12.075 ;
		RECT	14.765 12.175 14.815 12.305 ;
		RECT	14.765 9.755 14.815 9.885 ;
		RECT	19.685 12.175 19.735 12.305 ;
		RECT	19.685 9.755 19.735 9.885 ;
		RECT	14.965 12.175 15.015 12.305 ;
		RECT	14.965 9.755 15.015 9.885 ;
		RECT	19.485 12.175 19.535 12.305 ;
		RECT	19.485 9.755 19.535 9.885 ;
		RECT	14.565 9.065 14.615 9.195 ;
		RECT	19.885 9.065 19.935 9.195 ;
		RECT	14.765 9.295 14.815 9.425 ;
		RECT	14.765 6.875 14.815 7.005 ;
		RECT	19.685 9.295 19.735 9.425 ;
		RECT	19.685 6.875 19.735 7.005 ;
		RECT	14.965 9.295 15.015 9.425 ;
		RECT	14.965 6.875 15.015 7.005 ;
		RECT	19.485 9.295 19.535 9.425 ;
		RECT	19.485 6.875 19.535 7.005 ;
		RECT	14.565 6.185 14.615 6.315 ;
		RECT	19.885 6.185 19.935 6.315 ;
		RECT	14.765 6.415 14.815 6.545 ;
		RECT	14.765 3.995 14.815 4.125 ;
		RECT	19.685 6.415 19.735 6.545 ;
		RECT	19.685 3.995 19.735 4.125 ;
		RECT	14.965 6.415 15.015 6.545 ;
		RECT	14.965 3.995 15.015 4.125 ;
		RECT	19.485 6.415 19.535 6.545 ;
		RECT	19.485 3.995 19.535 4.125 ;
		RECT	14.565 164.585 14.615 164.715 ;
		RECT	19.885 164.585 19.935 164.715 ;
		RECT	14.765 164.815 14.815 164.945 ;
		RECT	14.765 162.395 14.815 162.525 ;
		RECT	19.685 164.815 19.735 164.945 ;
		RECT	19.685 162.395 19.735 162.525 ;
		RECT	14.965 164.815 15.015 164.945 ;
		RECT	14.965 162.395 15.015 162.525 ;
		RECT	19.485 164.815 19.535 164.945 ;
		RECT	19.485 162.395 19.535 162.525 ;
		RECT	14.565 161.705 14.615 161.835 ;
		RECT	19.885 161.705 19.935 161.835 ;
		RECT	14.765 161.935 14.815 162.065 ;
		RECT	14.765 159.515 14.815 159.645 ;
		RECT	19.685 161.935 19.735 162.065 ;
		RECT	19.685 159.515 19.735 159.645 ;
		RECT	14.965 161.935 15.015 162.065 ;
		RECT	14.965 159.515 15.015 159.645 ;
		RECT	19.485 161.935 19.535 162.065 ;
		RECT	19.485 159.515 19.535 159.645 ;
		RECT	14.565 158.825 14.615 158.955 ;
		RECT	19.885 158.825 19.935 158.955 ;
		RECT	14.765 159.055 14.815 159.185 ;
		RECT	14.765 156.635 14.815 156.765 ;
		RECT	19.685 159.055 19.735 159.185 ;
		RECT	19.685 156.635 19.735 156.765 ;
		RECT	14.965 159.055 15.015 159.185 ;
		RECT	14.965 156.635 15.015 156.765 ;
		RECT	19.485 159.055 19.535 159.185 ;
		RECT	19.485 156.635 19.535 156.765 ;
		RECT	20.085 182.095 20.265 182.225 ;
		RECT	20.875 181.865 21.055 181.995 ;
		RECT	20.085 179.675 20.265 179.805 ;
		RECT	20.43 179.445 20.48 179.575 ;
		RECT	20.085 156.175 20.265 156.305 ;
		RECT	20.875 155.945 21.055 156.075 ;
		RECT	20.085 153.755 20.265 153.885 ;
		RECT	20.43 153.525 20.48 153.655 ;
		RECT	20.085 153.295 20.265 153.425 ;
		RECT	20.875 153.065 21.055 153.195 ;
		RECT	20.085 150.875 20.265 151.005 ;
		RECT	20.43 150.645 20.48 150.775 ;
		RECT	20.085 150.415 20.265 150.545 ;
		RECT	20.875 150.185 21.055 150.315 ;
		RECT	20.085 147.995 20.265 148.125 ;
		RECT	20.43 147.765 20.48 147.895 ;
		RECT	20.085 147.535 20.265 147.665 ;
		RECT	20.875 147.305 21.055 147.435 ;
		RECT	20.085 145.115 20.265 145.245 ;
		RECT	20.43 144.885 20.48 145.015 ;
		RECT	20.085 144.655 20.265 144.785 ;
		RECT	20.875 144.425 21.055 144.555 ;
		RECT	20.085 142.235 20.265 142.365 ;
		RECT	20.43 142.005 20.48 142.135 ;
		RECT	20.085 141.775 20.265 141.905 ;
		RECT	20.875 141.545 21.055 141.675 ;
		RECT	20.085 139.355 20.265 139.485 ;
		RECT	20.43 139.125 20.48 139.255 ;
		RECT	20.085 138.895 20.265 139.025 ;
		RECT	20.875 138.665 21.055 138.795 ;
		RECT	20.085 136.475 20.265 136.605 ;
		RECT	20.43 136.245 20.48 136.375 ;
		RECT	20.085 136.015 20.265 136.145 ;
		RECT	20.875 135.785 21.055 135.915 ;
		RECT	20.085 133.595 20.265 133.725 ;
		RECT	20.43 133.365 20.48 133.495 ;
		RECT	20.085 133.135 20.265 133.265 ;
		RECT	20.875 132.905 21.055 133.035 ;
		RECT	20.085 130.715 20.265 130.845 ;
		RECT	20.43 130.485 20.48 130.615 ;
		RECT	20.085 130.255 20.265 130.385 ;
		RECT	20.875 130.025 21.055 130.155 ;
		RECT	20.085 127.835 20.265 127.965 ;
		RECT	20.43 127.605 20.48 127.735 ;
		RECT	20.085 179.215 20.265 179.345 ;
		RECT	20.875 178.985 21.055 179.115 ;
		RECT	20.085 176.795 20.265 176.925 ;
		RECT	20.43 176.565 20.48 176.695 ;
		RECT	20.085 127.375 20.265 127.505 ;
		RECT	20.875 127.145 21.055 127.275 ;
		RECT	20.085 124.955 20.265 125.085 ;
		RECT	20.43 124.725 20.48 124.855 ;
		RECT	20.085 124.495 20.265 124.625 ;
		RECT	20.875 124.265 21.055 124.395 ;
		RECT	20.085 122.075 20.265 122.205 ;
		RECT	20.43 121.845 20.48 121.975 ;
		RECT	20.085 121.615 20.265 121.745 ;
		RECT	20.875 121.385 21.055 121.515 ;
		RECT	20.085 119.195 20.265 119.325 ;
		RECT	20.43 118.965 20.48 119.095 ;
		RECT	20.085 118.735 20.265 118.865 ;
		RECT	20.875 118.505 21.055 118.635 ;
		RECT	20.085 116.315 20.265 116.445 ;
		RECT	20.43 116.085 20.48 116.215 ;
		RECT	20.085 115.855 20.265 115.985 ;
		RECT	20.875 115.625 21.055 115.755 ;
		RECT	20.085 113.435 20.265 113.565 ;
		RECT	20.43 113.205 20.48 113.335 ;
		RECT	20.085 112.975 20.265 113.105 ;
		RECT	20.875 112.745 21.055 112.875 ;
		RECT	20.085 110.555 20.265 110.685 ;
		RECT	20.43 110.325 20.48 110.455 ;
		RECT	20.085 110.095 20.265 110.225 ;
		RECT	20.875 109.865 21.055 109.995 ;
		RECT	20.085 107.675 20.265 107.805 ;
		RECT	20.43 107.445 20.48 107.575 ;
		RECT	20.085 107.215 20.265 107.345 ;
		RECT	20.875 106.985 21.055 107.115 ;
		RECT	20.085 104.795 20.265 104.925 ;
		RECT	20.43 104.565 20.48 104.695 ;
		RECT	20.085 104.335 20.265 104.465 ;
		RECT	20.875 104.105 21.055 104.235 ;
		RECT	20.085 101.915 20.265 102.045 ;
		RECT	20.43 101.685 20.48 101.815 ;
		RECT	20.085 101.455 20.265 101.585 ;
		RECT	20.875 101.225 21.055 101.355 ;
		RECT	20.085 99.035 20.265 99.165 ;
		RECT	20.43 98.805 20.48 98.935 ;
		RECT	20.085 176.335 20.265 176.465 ;
		RECT	20.875 176.105 21.055 176.235 ;
		RECT	20.085 173.915 20.265 174.045 ;
		RECT	20.43 173.685 20.48 173.815 ;
		RECT	20.085 98.575 20.265 98.705 ;
		RECT	20.875 98.345 21.055 98.475 ;
		RECT	20.085 96.155 20.265 96.285 ;
		RECT	20.43 95.925 20.48 96.055 ;
		RECT	20.085 95.695 20.265 95.825 ;
		RECT	20.875 95.465 21.055 95.595 ;
		RECT	20.085 93.275 20.265 93.405 ;
		RECT	20.43 93.045 20.48 93.175 ;
		RECT	20.085 92.815 20.265 92.945 ;
		RECT	20.875 92.585 21.055 92.715 ;
		RECT	20.085 90.395 20.265 90.525 ;
		RECT	20.43 90.165 20.48 90.295 ;
		RECT	20.085 89.935 20.265 90.065 ;
		RECT	20.875 89.705 21.055 89.835 ;
		RECT	20.085 87.515 20.265 87.645 ;
		RECT	20.43 87.285 20.48 87.415 ;
		RECT	20.085 87.055 20.265 87.185 ;
		RECT	20.875 86.825 21.055 86.955 ;
		RECT	20.085 84.635 20.265 84.765 ;
		RECT	20.43 84.405 20.48 84.535 ;
		RECT	20.085 84.175 20.265 84.305 ;
		RECT	20.875 83.945 21.055 84.075 ;
		RECT	20.085 81.755 20.265 81.885 ;
		RECT	20.43 81.525 20.48 81.655 ;
		RECT	20.085 81.295 20.265 81.425 ;
		RECT	20.875 81.065 21.055 81.195 ;
		RECT	20.085 78.875 20.265 79.005 ;
		RECT	20.43 78.645 20.48 78.775 ;
		RECT	20.085 78.415 20.265 78.545 ;
		RECT	20.875 78.185 21.055 78.315 ;
		RECT	20.085 75.995 20.265 76.125 ;
		RECT	20.43 75.765 20.48 75.895 ;
		RECT	20.085 75.535 20.265 75.665 ;
		RECT	20.875 75.305 21.055 75.435 ;
		RECT	20.085 73.115 20.265 73.245 ;
		RECT	20.43 72.885 20.48 73.015 ;
		RECT	20.085 72.655 20.265 72.785 ;
		RECT	20.875 72.425 21.055 72.555 ;
		RECT	20.085 70.235 20.265 70.365 ;
		RECT	20.43 70.005 20.48 70.135 ;
		RECT	20.085 173.455 20.265 173.585 ;
		RECT	20.875 173.225 21.055 173.355 ;
		RECT	20.085 171.035 20.265 171.165 ;
		RECT	20.43 170.805 20.48 170.935 ;
		RECT	20.085 69.775 20.265 69.905 ;
		RECT	20.875 69.545 21.055 69.675 ;
		RECT	20.085 67.355 20.265 67.485 ;
		RECT	20.43 67.125 20.48 67.255 ;
		RECT	20.085 66.895 20.265 67.025 ;
		RECT	20.875 66.665 21.055 66.795 ;
		RECT	20.085 64.475 20.265 64.605 ;
		RECT	20.43 64.245 20.48 64.375 ;
		RECT	20.085 64.015 20.265 64.145 ;
		RECT	20.875 63.785 21.055 63.915 ;
		RECT	20.085 61.595 20.265 61.725 ;
		RECT	20.43 61.365 20.48 61.495 ;
		RECT	20.085 61.135 20.265 61.265 ;
		RECT	20.875 60.905 21.055 61.035 ;
		RECT	20.085 58.715 20.265 58.845 ;
		RECT	20.43 58.485 20.48 58.615 ;
		RECT	20.085 58.255 20.265 58.385 ;
		RECT	20.875 58.025 21.055 58.155 ;
		RECT	20.085 55.835 20.265 55.965 ;
		RECT	20.43 55.605 20.48 55.735 ;
		RECT	20.085 55.375 20.265 55.505 ;
		RECT	20.875 55.145 21.055 55.275 ;
		RECT	20.085 52.955 20.265 53.085 ;
		RECT	20.43 52.725 20.48 52.855 ;
		RECT	20.085 52.495 20.265 52.625 ;
		RECT	20.875 52.265 21.055 52.395 ;
		RECT	20.085 50.075 20.265 50.205 ;
		RECT	20.43 49.845 20.48 49.975 ;
		RECT	20.085 49.615 20.265 49.745 ;
		RECT	20.875 49.385 21.055 49.515 ;
		RECT	20.085 47.195 20.265 47.325 ;
		RECT	20.43 46.965 20.48 47.095 ;
		RECT	20.085 46.735 20.265 46.865 ;
		RECT	20.875 46.505 21.055 46.635 ;
		RECT	20.085 44.315 20.265 44.445 ;
		RECT	20.43 44.085 20.48 44.215 ;
		RECT	20.085 43.855 20.265 43.985 ;
		RECT	20.875 43.625 21.055 43.755 ;
		RECT	20.085 41.435 20.265 41.565 ;
		RECT	20.43 41.205 20.48 41.335 ;
		RECT	20.085 170.575 20.265 170.705 ;
		RECT	20.875 170.345 21.055 170.475 ;
		RECT	20.085 168.155 20.265 168.285 ;
		RECT	20.43 167.925 20.48 168.055 ;
		RECT	20.085 40.975 20.265 41.105 ;
		RECT	20.875 40.745 21.055 40.875 ;
		RECT	20.085 38.555 20.265 38.685 ;
		RECT	20.43 38.325 20.48 38.455 ;
		RECT	20.085 38.095 20.265 38.225 ;
		RECT	20.875 37.865 21.055 37.995 ;
		RECT	20.085 35.675 20.265 35.805 ;
		RECT	20.43 35.445 20.48 35.575 ;
		RECT	20.085 35.215 20.265 35.345 ;
		RECT	20.875 34.985 21.055 35.115 ;
		RECT	20.085 32.795 20.265 32.925 ;
		RECT	20.43 32.565 20.48 32.695 ;
		RECT	20.085 32.335 20.265 32.465 ;
		RECT	20.875 32.105 21.055 32.235 ;
		RECT	20.085 29.915 20.265 30.045 ;
		RECT	20.43 29.685 20.48 29.815 ;
		RECT	20.085 29.455 20.265 29.585 ;
		RECT	20.875 29.225 21.055 29.355 ;
		RECT	20.085 27.035 20.265 27.165 ;
		RECT	20.43 26.805 20.48 26.935 ;
		RECT	20.085 26.575 20.265 26.705 ;
		RECT	20.875 26.345 21.055 26.475 ;
		RECT	20.085 24.155 20.265 24.285 ;
		RECT	20.43 23.925 20.48 24.055 ;
		RECT	20.085 23.695 20.265 23.825 ;
		RECT	20.875 23.465 21.055 23.595 ;
		RECT	20.085 21.275 20.265 21.405 ;
		RECT	20.43 21.045 20.48 21.175 ;
		RECT	20.085 20.815 20.265 20.945 ;
		RECT	20.875 20.585 21.055 20.715 ;
		RECT	20.085 18.395 20.265 18.525 ;
		RECT	20.43 18.165 20.48 18.295 ;
		RECT	20.085 17.935 20.265 18.065 ;
		RECT	20.875 17.705 21.055 17.835 ;
		RECT	20.085 15.515 20.265 15.645 ;
		RECT	20.43 15.285 20.48 15.415 ;
		RECT	20.085 15.055 20.265 15.185 ;
		RECT	20.875 14.825 21.055 14.955 ;
		RECT	20.085 12.635 20.265 12.765 ;
		RECT	20.43 12.405 20.48 12.535 ;
		RECT	20.085 167.695 20.265 167.825 ;
		RECT	20.875 167.465 21.055 167.595 ;
		RECT	20.085 165.275 20.265 165.405 ;
		RECT	20.43 165.045 20.48 165.175 ;
		RECT	20.085 12.175 20.265 12.305 ;
		RECT	20.875 11.945 21.055 12.075 ;
		RECT	20.085 9.755 20.265 9.885 ;
		RECT	20.43 9.525 20.48 9.655 ;
		RECT	20.085 9.295 20.265 9.425 ;
		RECT	20.875 9.065 21.055 9.195 ;
		RECT	20.085 6.875 20.265 7.005 ;
		RECT	20.43 6.645 20.48 6.775 ;
		RECT	20.085 6.415 20.265 6.545 ;
		RECT	20.875 6.185 21.055 6.315 ;
		RECT	20.085 3.995 20.265 4.125 ;
		RECT	20.43 3.765 20.48 3.895 ;
		RECT	20.085 164.815 20.265 164.945 ;
		RECT	20.875 164.585 21.055 164.715 ;
		RECT	20.085 162.395 20.265 162.525 ;
		RECT	20.43 162.165 20.48 162.295 ;
		RECT	20.085 161.935 20.265 162.065 ;
		RECT	20.875 161.705 21.055 161.835 ;
		RECT	20.085 159.515 20.265 159.645 ;
		RECT	20.43 159.285 20.48 159.415 ;
		RECT	20.085 159.055 20.265 159.185 ;
		RECT	20.875 158.825 21.055 158.955 ;
		RECT	20.085 156.635 20.265 156.765 ;
		RECT	20.43 156.405 20.48 156.535 ;
		RECT	20.085 3.535 20.265 3.665 ;
		RECT	20.875 3.305 21.055 3.435 ;
		RECT	20.085 1.115 20.265 1.245 ;
		RECT	20.43 0.885 20.48 1.015 ;
		RECT	20.085 184.975 20.265 185.105 ;
		RECT	20.875 184.745 21.055 184.875 ;
		RECT	20.085 182.555 20.265 182.685 ;
		RECT	20.43 182.325 20.48 182.455 ;
		RECT	14.565 411.425 14.615 411.555 ;
		RECT	19.885 411.425 19.935 411.555 ;
		RECT	14.765 411.195 14.815 411.325 ;
		RECT	14.765 413.615 14.815 413.745 ;
		RECT	19.685 411.195 19.735 411.325 ;
		RECT	19.685 413.615 19.735 413.745 ;
		RECT	14.965 411.195 15.015 411.325 ;
		RECT	14.965 413.615 15.015 413.745 ;
		RECT	19.485 411.195 19.535 411.325 ;
		RECT	19.485 413.615 19.535 413.745 ;
		RECT	14.565 229.985 14.615 230.115 ;
		RECT	19.885 229.985 19.935 230.115 ;
		RECT	14.765 229.755 14.815 229.885 ;
		RECT	14.765 232.175 14.815 232.305 ;
		RECT	19.685 229.755 19.735 229.885 ;
		RECT	19.685 232.175 19.735 232.305 ;
		RECT	14.965 229.755 15.015 229.885 ;
		RECT	14.965 232.175 15.015 232.305 ;
		RECT	19.485 229.755 19.535 229.885 ;
		RECT	19.485 232.175 19.535 232.305 ;
		RECT	14.565 232.865 14.615 232.995 ;
		RECT	19.885 232.865 19.935 232.995 ;
		RECT	14.765 232.635 14.815 232.765 ;
		RECT	14.765 235.055 14.815 235.185 ;
		RECT	19.685 232.635 19.735 232.765 ;
		RECT	19.685 235.055 19.735 235.185 ;
		RECT	14.965 232.635 15.015 232.765 ;
		RECT	14.965 235.055 15.015 235.185 ;
		RECT	19.485 232.635 19.535 232.765 ;
		RECT	19.485 235.055 19.535 235.185 ;
		RECT	14.565 258.785 14.615 258.915 ;
		RECT	19.885 258.785 19.935 258.915 ;
		RECT	14.765 258.555 14.815 258.685 ;
		RECT	14.765 260.975 14.815 261.105 ;
		RECT	19.685 258.555 19.735 258.685 ;
		RECT	19.685 260.975 19.735 261.105 ;
		RECT	14.965 258.555 15.015 258.685 ;
		RECT	14.965 260.975 15.015 261.105 ;
		RECT	19.485 258.555 19.535 258.685 ;
		RECT	19.485 260.975 19.535 261.105 ;
		RECT	14.565 261.665 14.615 261.795 ;
		RECT	19.885 261.665 19.935 261.795 ;
		RECT	14.765 261.435 14.815 261.565 ;
		RECT	14.765 263.855 14.815 263.985 ;
		RECT	19.685 261.435 19.735 261.565 ;
		RECT	19.685 263.855 19.735 263.985 ;
		RECT	14.965 261.435 15.015 261.565 ;
		RECT	14.965 263.855 15.015 263.985 ;
		RECT	19.485 261.435 19.535 261.565 ;
		RECT	19.485 263.855 19.535 263.985 ;
		RECT	14.565 264.545 14.615 264.675 ;
		RECT	19.885 264.545 19.935 264.675 ;
		RECT	14.765 264.315 14.815 264.445 ;
		RECT	14.765 266.735 14.815 266.865 ;
		RECT	19.685 264.315 19.735 264.445 ;
		RECT	19.685 266.735 19.735 266.865 ;
		RECT	14.965 264.315 15.015 264.445 ;
		RECT	14.965 266.735 15.015 266.865 ;
		RECT	19.485 264.315 19.535 264.445 ;
		RECT	19.485 266.735 19.535 266.865 ;
		RECT	14.565 267.425 14.615 267.555 ;
		RECT	19.885 267.425 19.935 267.555 ;
		RECT	14.765 267.195 14.815 267.325 ;
		RECT	14.765 269.615 14.815 269.745 ;
		RECT	19.685 267.195 19.735 267.325 ;
		RECT	19.685 269.615 19.735 269.745 ;
		RECT	14.965 267.195 15.015 267.325 ;
		RECT	14.965 269.615 15.015 269.745 ;
		RECT	19.485 267.195 19.535 267.325 ;
		RECT	19.485 269.615 19.535 269.745 ;
		RECT	14.565 270.305 14.615 270.435 ;
		RECT	19.885 270.305 19.935 270.435 ;
		RECT	14.765 270.075 14.815 270.205 ;
		RECT	14.765 272.495 14.815 272.625 ;
		RECT	19.685 270.075 19.735 270.205 ;
		RECT	19.685 272.495 19.735 272.625 ;
		RECT	14.965 270.075 15.015 270.205 ;
		RECT	14.965 272.495 15.015 272.625 ;
		RECT	19.485 270.075 19.535 270.205 ;
		RECT	19.485 272.495 19.535 272.625 ;
		RECT	14.565 273.185 14.615 273.315 ;
		RECT	19.885 273.185 19.935 273.315 ;
		RECT	14.765 272.955 14.815 273.085 ;
		RECT	14.765 275.375 14.815 275.505 ;
		RECT	19.685 272.955 19.735 273.085 ;
		RECT	19.685 275.375 19.735 275.505 ;
		RECT	14.965 272.955 15.015 273.085 ;
		RECT	14.965 275.375 15.015 275.505 ;
		RECT	19.485 272.955 19.535 273.085 ;
		RECT	19.485 275.375 19.535 275.505 ;
		RECT	14.565 276.065 14.615 276.195 ;
		RECT	19.885 276.065 19.935 276.195 ;
		RECT	14.765 275.835 14.815 275.965 ;
		RECT	14.765 278.255 14.815 278.385 ;
		RECT	19.685 275.835 19.735 275.965 ;
		RECT	19.685 278.255 19.735 278.385 ;
		RECT	14.965 275.835 15.015 275.965 ;
		RECT	14.965 278.255 15.015 278.385 ;
		RECT	19.485 275.835 19.535 275.965 ;
		RECT	19.485 278.255 19.535 278.385 ;
		RECT	14.565 278.945 14.615 279.075 ;
		RECT	19.885 278.945 19.935 279.075 ;
		RECT	14.765 278.715 14.815 278.845 ;
		RECT	14.765 281.135 14.815 281.265 ;
		RECT	19.685 278.715 19.735 278.845 ;
		RECT	19.685 281.135 19.735 281.265 ;
		RECT	14.965 278.715 15.015 278.845 ;
		RECT	14.965 281.135 15.015 281.265 ;
		RECT	19.485 278.715 19.535 278.845 ;
		RECT	19.485 281.135 19.535 281.265 ;
		RECT	14.565 281.825 14.615 281.955 ;
		RECT	19.885 281.825 19.935 281.955 ;
		RECT	14.765 281.595 14.815 281.725 ;
		RECT	14.765 284.015 14.815 284.145 ;
		RECT	19.685 281.595 19.735 281.725 ;
		RECT	19.685 284.015 19.735 284.145 ;
		RECT	14.965 281.595 15.015 281.725 ;
		RECT	14.965 284.015 15.015 284.145 ;
		RECT	19.485 281.595 19.535 281.725 ;
		RECT	19.485 284.015 19.535 284.145 ;
		RECT	14.565 284.705 14.615 284.835 ;
		RECT	19.885 284.705 19.935 284.835 ;
		RECT	14.765 284.475 14.815 284.605 ;
		RECT	14.765 286.895 14.815 287.025 ;
		RECT	19.685 284.475 19.735 284.605 ;
		RECT	19.685 286.895 19.735 287.025 ;
		RECT	14.965 284.475 15.015 284.605 ;
		RECT	14.965 286.895 15.015 287.025 ;
		RECT	19.485 284.475 19.535 284.605 ;
		RECT	19.485 286.895 19.535 287.025 ;
		RECT	14.565 235.745 14.615 235.875 ;
		RECT	19.885 235.745 19.935 235.875 ;
		RECT	14.765 235.515 14.815 235.645 ;
		RECT	14.765 237.935 14.815 238.065 ;
		RECT	19.685 235.515 19.735 235.645 ;
		RECT	19.685 237.935 19.735 238.065 ;
		RECT	14.965 235.515 15.015 235.645 ;
		RECT	14.965 237.935 15.015 238.065 ;
		RECT	19.485 235.515 19.535 235.645 ;
		RECT	19.485 237.935 19.535 238.065 ;
		RECT	14.565 287.585 14.615 287.715 ;
		RECT	19.885 287.585 19.935 287.715 ;
		RECT	14.765 287.355 14.815 287.485 ;
		RECT	14.765 289.775 14.815 289.905 ;
		RECT	19.685 287.355 19.735 287.485 ;
		RECT	19.685 289.775 19.735 289.905 ;
		RECT	14.965 287.355 15.015 287.485 ;
		RECT	14.965 289.775 15.015 289.905 ;
		RECT	19.485 287.355 19.535 287.485 ;
		RECT	19.485 289.775 19.535 289.905 ;
		RECT	14.565 290.465 14.615 290.595 ;
		RECT	19.885 290.465 19.935 290.595 ;
		RECT	14.765 290.235 14.815 290.365 ;
		RECT	14.765 292.655 14.815 292.785 ;
		RECT	19.685 290.235 19.735 290.365 ;
		RECT	19.685 292.655 19.735 292.785 ;
		RECT	14.965 290.235 15.015 290.365 ;
		RECT	14.965 292.655 15.015 292.785 ;
		RECT	19.485 290.235 19.535 290.365 ;
		RECT	19.485 292.655 19.535 292.785 ;
		RECT	14.565 293.345 14.615 293.475 ;
		RECT	19.885 293.345 19.935 293.475 ;
		RECT	14.765 293.115 14.815 293.245 ;
		RECT	14.765 295.535 14.815 295.665 ;
		RECT	19.685 293.115 19.735 293.245 ;
		RECT	19.685 295.535 19.735 295.665 ;
		RECT	14.965 293.115 15.015 293.245 ;
		RECT	14.965 295.535 15.015 295.665 ;
		RECT	19.485 293.115 19.535 293.245 ;
		RECT	19.485 295.535 19.535 295.665 ;
		RECT	14.565 296.225 14.615 296.355 ;
		RECT	19.885 296.225 19.935 296.355 ;
		RECT	14.765 295.995 14.815 296.125 ;
		RECT	14.765 298.415 14.815 298.545 ;
		RECT	19.685 295.995 19.735 296.125 ;
		RECT	19.685 298.415 19.735 298.545 ;
		RECT	14.965 295.995 15.015 296.125 ;
		RECT	14.965 298.415 15.015 298.545 ;
		RECT	19.485 295.995 19.535 296.125 ;
		RECT	19.485 298.415 19.535 298.545 ;
		RECT	14.565 299.105 14.615 299.235 ;
		RECT	19.885 299.105 19.935 299.235 ;
		RECT	14.765 298.875 14.815 299.005 ;
		RECT	14.765 301.295 14.815 301.425 ;
		RECT	19.685 298.875 19.735 299.005 ;
		RECT	19.685 301.295 19.735 301.425 ;
		RECT	14.965 298.875 15.015 299.005 ;
		RECT	14.965 301.295 15.015 301.425 ;
		RECT	19.485 298.875 19.535 299.005 ;
		RECT	19.485 301.295 19.535 301.425 ;
		RECT	14.565 301.985 14.615 302.115 ;
		RECT	19.885 301.985 19.935 302.115 ;
		RECT	14.765 301.755 14.815 301.885 ;
		RECT	14.765 304.175 14.815 304.305 ;
		RECT	19.685 301.755 19.735 301.885 ;
		RECT	19.685 304.175 19.735 304.305 ;
		RECT	14.965 301.755 15.015 301.885 ;
		RECT	14.965 304.175 15.015 304.305 ;
		RECT	19.485 301.755 19.535 301.885 ;
		RECT	19.485 304.175 19.535 304.305 ;
		RECT	14.565 304.865 14.615 304.995 ;
		RECT	19.885 304.865 19.935 304.995 ;
		RECT	14.765 304.635 14.815 304.765 ;
		RECT	14.765 307.055 14.815 307.185 ;
		RECT	19.685 304.635 19.735 304.765 ;
		RECT	19.685 307.055 19.735 307.185 ;
		RECT	14.965 304.635 15.015 304.765 ;
		RECT	14.965 307.055 15.015 307.185 ;
		RECT	19.485 304.635 19.535 304.765 ;
		RECT	19.485 307.055 19.535 307.185 ;
		RECT	14.565 307.745 14.615 307.875 ;
		RECT	19.885 307.745 19.935 307.875 ;
		RECT	14.765 307.515 14.815 307.645 ;
		RECT	14.765 309.935 14.815 310.065 ;
		RECT	19.685 307.515 19.735 307.645 ;
		RECT	19.685 309.935 19.735 310.065 ;
		RECT	14.965 307.515 15.015 307.645 ;
		RECT	14.965 309.935 15.015 310.065 ;
		RECT	19.485 307.515 19.535 307.645 ;
		RECT	19.485 309.935 19.535 310.065 ;
		RECT	14.565 310.625 14.615 310.755 ;
		RECT	19.885 310.625 19.935 310.755 ;
		RECT	14.765 310.395 14.815 310.525 ;
		RECT	14.765 312.815 14.815 312.945 ;
		RECT	19.685 310.395 19.735 310.525 ;
		RECT	19.685 312.815 19.735 312.945 ;
		RECT	14.965 310.395 15.015 310.525 ;
		RECT	14.965 312.815 15.015 312.945 ;
		RECT	19.485 310.395 19.535 310.525 ;
		RECT	19.485 312.815 19.535 312.945 ;
		RECT	14.565 313.505 14.615 313.635 ;
		RECT	19.885 313.505 19.935 313.635 ;
		RECT	14.765 313.275 14.815 313.405 ;
		RECT	14.765 315.695 14.815 315.825 ;
		RECT	19.685 313.275 19.735 313.405 ;
		RECT	19.685 315.695 19.735 315.825 ;
		RECT	14.965 313.275 15.015 313.405 ;
		RECT	14.965 315.695 15.015 315.825 ;
		RECT	19.485 313.275 19.535 313.405 ;
		RECT	19.485 315.695 19.535 315.825 ;
		RECT	14.565 238.625 14.615 238.755 ;
		RECT	19.885 238.625 19.935 238.755 ;
		RECT	14.765 238.395 14.815 238.525 ;
		RECT	14.765 240.815 14.815 240.945 ;
		RECT	19.685 238.395 19.735 238.525 ;
		RECT	19.685 240.815 19.735 240.945 ;
		RECT	14.965 238.395 15.015 238.525 ;
		RECT	14.965 240.815 15.015 240.945 ;
		RECT	19.485 238.395 19.535 238.525 ;
		RECT	19.485 240.815 19.535 240.945 ;
		RECT	14.565 316.385 14.615 316.515 ;
		RECT	19.885 316.385 19.935 316.515 ;
		RECT	14.765 316.155 14.815 316.285 ;
		RECT	14.765 318.575 14.815 318.705 ;
		RECT	19.685 316.155 19.735 316.285 ;
		RECT	19.685 318.575 19.735 318.705 ;
		RECT	14.965 316.155 15.015 316.285 ;
		RECT	14.965 318.575 15.015 318.705 ;
		RECT	19.485 316.155 19.535 316.285 ;
		RECT	19.485 318.575 19.535 318.705 ;
		RECT	14.565 319.265 14.615 319.395 ;
		RECT	19.885 319.265 19.935 319.395 ;
		RECT	14.765 319.035 14.815 319.165 ;
		RECT	14.765 321.455 14.815 321.585 ;
		RECT	19.685 319.035 19.735 319.165 ;
		RECT	19.685 321.455 19.735 321.585 ;
		RECT	14.965 319.035 15.015 319.165 ;
		RECT	14.965 321.455 15.015 321.585 ;
		RECT	19.485 319.035 19.535 319.165 ;
		RECT	19.485 321.455 19.535 321.585 ;
		RECT	14.565 322.145 14.615 322.275 ;
		RECT	19.885 322.145 19.935 322.275 ;
		RECT	14.765 321.915 14.815 322.045 ;
		RECT	14.765 324.335 14.815 324.465 ;
		RECT	19.685 321.915 19.735 322.045 ;
		RECT	19.685 324.335 19.735 324.465 ;
		RECT	14.965 321.915 15.015 322.045 ;
		RECT	14.965 324.335 15.015 324.465 ;
		RECT	19.485 321.915 19.535 322.045 ;
		RECT	19.485 324.335 19.535 324.465 ;
		RECT	14.565 325.025 14.615 325.155 ;
		RECT	19.885 325.025 19.935 325.155 ;
		RECT	14.765 324.795 14.815 324.925 ;
		RECT	14.765 327.215 14.815 327.345 ;
		RECT	19.685 324.795 19.735 324.925 ;
		RECT	19.685 327.215 19.735 327.345 ;
		RECT	14.965 324.795 15.015 324.925 ;
		RECT	14.965 327.215 15.015 327.345 ;
		RECT	19.485 324.795 19.535 324.925 ;
		RECT	19.485 327.215 19.535 327.345 ;
		RECT	14.565 327.905 14.615 328.035 ;
		RECT	19.885 327.905 19.935 328.035 ;
		RECT	14.765 327.675 14.815 327.805 ;
		RECT	14.765 330.095 14.815 330.225 ;
		RECT	19.685 327.675 19.735 327.805 ;
		RECT	19.685 330.095 19.735 330.225 ;
		RECT	14.965 327.675 15.015 327.805 ;
		RECT	14.965 330.095 15.015 330.225 ;
		RECT	19.485 327.675 19.535 327.805 ;
		RECT	19.485 330.095 19.535 330.225 ;
		RECT	14.565 330.785 14.615 330.915 ;
		RECT	19.885 330.785 19.935 330.915 ;
		RECT	14.765 330.555 14.815 330.685 ;
		RECT	14.765 332.975 14.815 333.105 ;
		RECT	19.685 330.555 19.735 330.685 ;
		RECT	19.685 332.975 19.735 333.105 ;
		RECT	14.965 330.555 15.015 330.685 ;
		RECT	14.965 332.975 15.015 333.105 ;
		RECT	19.485 330.555 19.535 330.685 ;
		RECT	19.485 332.975 19.535 333.105 ;
		RECT	14.565 333.665 14.615 333.795 ;
		RECT	19.885 333.665 19.935 333.795 ;
		RECT	14.765 333.435 14.815 333.565 ;
		RECT	14.765 335.855 14.815 335.985 ;
		RECT	19.685 333.435 19.735 333.565 ;
		RECT	19.685 335.855 19.735 335.985 ;
		RECT	14.965 333.435 15.015 333.565 ;
		RECT	14.965 335.855 15.015 335.985 ;
		RECT	19.485 333.435 19.535 333.565 ;
		RECT	19.485 335.855 19.535 335.985 ;
		RECT	14.565 336.545 14.615 336.675 ;
		RECT	19.885 336.545 19.935 336.675 ;
		RECT	14.765 336.315 14.815 336.445 ;
		RECT	14.765 338.735 14.815 338.865 ;
		RECT	19.685 336.315 19.735 336.445 ;
		RECT	19.685 338.735 19.735 338.865 ;
		RECT	14.965 336.315 15.015 336.445 ;
		RECT	14.965 338.735 15.015 338.865 ;
		RECT	19.485 336.315 19.535 336.445 ;
		RECT	19.485 338.735 19.535 338.865 ;
		RECT	14.565 339.425 14.615 339.555 ;
		RECT	19.885 339.425 19.935 339.555 ;
		RECT	14.765 339.195 14.815 339.325 ;
		RECT	14.765 341.615 14.815 341.745 ;
		RECT	19.685 339.195 19.735 339.325 ;
		RECT	19.685 341.615 19.735 341.745 ;
		RECT	14.965 339.195 15.015 339.325 ;
		RECT	14.965 341.615 15.015 341.745 ;
		RECT	19.485 339.195 19.535 339.325 ;
		RECT	19.485 341.615 19.535 341.745 ;
		RECT	14.565 342.305 14.615 342.435 ;
		RECT	19.885 342.305 19.935 342.435 ;
		RECT	14.765 342.075 14.815 342.205 ;
		RECT	14.765 344.495 14.815 344.625 ;
		RECT	19.685 342.075 19.735 342.205 ;
		RECT	19.685 344.495 19.735 344.625 ;
		RECT	14.965 342.075 15.015 342.205 ;
		RECT	14.965 344.495 15.015 344.625 ;
		RECT	19.485 342.075 19.535 342.205 ;
		RECT	19.485 344.495 19.535 344.625 ;
		RECT	14.565 241.505 14.615 241.635 ;
		RECT	19.885 241.505 19.935 241.635 ;
		RECT	14.765 241.275 14.815 241.405 ;
		RECT	14.765 243.695 14.815 243.825 ;
		RECT	19.685 241.275 19.735 241.405 ;
		RECT	19.685 243.695 19.735 243.825 ;
		RECT	14.965 241.275 15.015 241.405 ;
		RECT	14.965 243.695 15.015 243.825 ;
		RECT	19.485 241.275 19.535 241.405 ;
		RECT	19.485 243.695 19.535 243.825 ;
		RECT	14.565 345.185 14.615 345.315 ;
		RECT	19.885 345.185 19.935 345.315 ;
		RECT	14.765 344.955 14.815 345.085 ;
		RECT	14.765 347.375 14.815 347.505 ;
		RECT	19.685 344.955 19.735 345.085 ;
		RECT	19.685 347.375 19.735 347.505 ;
		RECT	14.965 344.955 15.015 345.085 ;
		RECT	14.965 347.375 15.015 347.505 ;
		RECT	19.485 344.955 19.535 345.085 ;
		RECT	19.485 347.375 19.535 347.505 ;
		RECT	14.565 348.065 14.615 348.195 ;
		RECT	19.885 348.065 19.935 348.195 ;
		RECT	14.765 347.835 14.815 347.965 ;
		RECT	14.765 350.255 14.815 350.385 ;
		RECT	19.685 347.835 19.735 347.965 ;
		RECT	19.685 350.255 19.735 350.385 ;
		RECT	14.965 347.835 15.015 347.965 ;
		RECT	14.965 350.255 15.015 350.385 ;
		RECT	19.485 347.835 19.535 347.965 ;
		RECT	19.485 350.255 19.535 350.385 ;
		RECT	14.565 350.945 14.615 351.075 ;
		RECT	19.885 350.945 19.935 351.075 ;
		RECT	14.765 350.715 14.815 350.845 ;
		RECT	14.765 353.135 14.815 353.265 ;
		RECT	19.685 350.715 19.735 350.845 ;
		RECT	19.685 353.135 19.735 353.265 ;
		RECT	14.965 350.715 15.015 350.845 ;
		RECT	14.965 353.135 15.015 353.265 ;
		RECT	19.485 350.715 19.535 350.845 ;
		RECT	19.485 353.135 19.535 353.265 ;
		RECT	14.565 353.825 14.615 353.955 ;
		RECT	19.885 353.825 19.935 353.955 ;
		RECT	14.765 353.595 14.815 353.725 ;
		RECT	14.765 356.015 14.815 356.145 ;
		RECT	19.685 353.595 19.735 353.725 ;
		RECT	19.685 356.015 19.735 356.145 ;
		RECT	14.965 353.595 15.015 353.725 ;
		RECT	14.965 356.015 15.015 356.145 ;
		RECT	19.485 353.595 19.535 353.725 ;
		RECT	19.485 356.015 19.535 356.145 ;
		RECT	14.565 356.705 14.615 356.835 ;
		RECT	19.885 356.705 19.935 356.835 ;
		RECT	14.765 356.475 14.815 356.605 ;
		RECT	14.765 358.895 14.815 359.025 ;
		RECT	19.685 356.475 19.735 356.605 ;
		RECT	19.685 358.895 19.735 359.025 ;
		RECT	14.965 356.475 15.015 356.605 ;
		RECT	14.965 358.895 15.015 359.025 ;
		RECT	19.485 356.475 19.535 356.605 ;
		RECT	19.485 358.895 19.535 359.025 ;
		RECT	14.565 359.585 14.615 359.715 ;
		RECT	19.885 359.585 19.935 359.715 ;
		RECT	14.765 359.355 14.815 359.485 ;
		RECT	14.765 361.775 14.815 361.905 ;
		RECT	19.685 359.355 19.735 359.485 ;
		RECT	19.685 361.775 19.735 361.905 ;
		RECT	14.965 359.355 15.015 359.485 ;
		RECT	14.965 361.775 15.015 361.905 ;
		RECT	19.485 359.355 19.535 359.485 ;
		RECT	19.485 361.775 19.535 361.905 ;
		RECT	14.565 362.465 14.615 362.595 ;
		RECT	19.885 362.465 19.935 362.595 ;
		RECT	14.765 362.235 14.815 362.365 ;
		RECT	14.765 364.655 14.815 364.785 ;
		RECT	19.685 362.235 19.735 362.365 ;
		RECT	19.685 364.655 19.735 364.785 ;
		RECT	14.965 362.235 15.015 362.365 ;
		RECT	14.965 364.655 15.015 364.785 ;
		RECT	19.485 362.235 19.535 362.365 ;
		RECT	19.485 364.655 19.535 364.785 ;
		RECT	14.565 365.345 14.615 365.475 ;
		RECT	19.885 365.345 19.935 365.475 ;
		RECT	14.765 365.115 14.815 365.245 ;
		RECT	14.765 367.535 14.815 367.665 ;
		RECT	19.685 365.115 19.735 365.245 ;
		RECT	19.685 367.535 19.735 367.665 ;
		RECT	14.965 365.115 15.015 365.245 ;
		RECT	14.965 367.535 15.015 367.665 ;
		RECT	19.485 365.115 19.535 365.245 ;
		RECT	19.485 367.535 19.535 367.665 ;
		RECT	14.565 368.225 14.615 368.355 ;
		RECT	19.885 368.225 19.935 368.355 ;
		RECT	14.765 367.995 14.815 368.125 ;
		RECT	14.765 370.415 14.815 370.545 ;
		RECT	19.685 367.995 19.735 368.125 ;
		RECT	19.685 370.415 19.735 370.545 ;
		RECT	14.965 367.995 15.015 368.125 ;
		RECT	14.965 370.415 15.015 370.545 ;
		RECT	19.485 367.995 19.535 368.125 ;
		RECT	19.485 370.415 19.535 370.545 ;
		RECT	14.565 371.105 14.615 371.235 ;
		RECT	19.885 371.105 19.935 371.235 ;
		RECT	14.765 370.875 14.815 371.005 ;
		RECT	14.765 373.295 14.815 373.425 ;
		RECT	19.685 370.875 19.735 371.005 ;
		RECT	19.685 373.295 19.735 373.425 ;
		RECT	14.965 370.875 15.015 371.005 ;
		RECT	14.965 373.295 15.015 373.425 ;
		RECT	19.485 370.875 19.535 371.005 ;
		RECT	19.485 373.295 19.535 373.425 ;
		RECT	14.565 244.385 14.615 244.515 ;
		RECT	19.885 244.385 19.935 244.515 ;
		RECT	14.765 244.155 14.815 244.285 ;
		RECT	14.765 246.575 14.815 246.705 ;
		RECT	19.685 244.155 19.735 244.285 ;
		RECT	19.685 246.575 19.735 246.705 ;
		RECT	14.965 244.155 15.015 244.285 ;
		RECT	14.965 246.575 15.015 246.705 ;
		RECT	19.485 244.155 19.535 244.285 ;
		RECT	19.485 246.575 19.535 246.705 ;
		RECT	14.565 373.985 14.615 374.115 ;
		RECT	19.885 373.985 19.935 374.115 ;
		RECT	14.765 373.755 14.815 373.885 ;
		RECT	14.765 376.175 14.815 376.305 ;
		RECT	19.685 373.755 19.735 373.885 ;
		RECT	19.685 376.175 19.735 376.305 ;
		RECT	14.965 373.755 15.015 373.885 ;
		RECT	14.965 376.175 15.015 376.305 ;
		RECT	19.485 373.755 19.535 373.885 ;
		RECT	19.485 376.175 19.535 376.305 ;
		RECT	14.565 376.865 14.615 376.995 ;
		RECT	19.885 376.865 19.935 376.995 ;
		RECT	14.765 376.635 14.815 376.765 ;
		RECT	14.765 379.055 14.815 379.185 ;
		RECT	19.685 376.635 19.735 376.765 ;
		RECT	19.685 379.055 19.735 379.185 ;
		RECT	14.965 376.635 15.015 376.765 ;
		RECT	14.965 379.055 15.015 379.185 ;
		RECT	19.485 376.635 19.535 376.765 ;
		RECT	19.485 379.055 19.535 379.185 ;
		RECT	14.565 379.745 14.615 379.875 ;
		RECT	19.885 379.745 19.935 379.875 ;
		RECT	14.765 379.515 14.815 379.645 ;
		RECT	14.765 381.935 14.815 382.065 ;
		RECT	19.685 379.515 19.735 379.645 ;
		RECT	19.685 381.935 19.735 382.065 ;
		RECT	14.965 379.515 15.015 379.645 ;
		RECT	14.965 381.935 15.015 382.065 ;
		RECT	19.485 379.515 19.535 379.645 ;
		RECT	19.485 381.935 19.535 382.065 ;
		RECT	14.565 382.625 14.615 382.755 ;
		RECT	19.885 382.625 19.935 382.755 ;
		RECT	14.765 382.395 14.815 382.525 ;
		RECT	14.765 384.815 14.815 384.945 ;
		RECT	19.685 382.395 19.735 382.525 ;
		RECT	19.685 384.815 19.735 384.945 ;
		RECT	14.965 382.395 15.015 382.525 ;
		RECT	14.965 384.815 15.015 384.945 ;
		RECT	19.485 382.395 19.535 382.525 ;
		RECT	19.485 384.815 19.535 384.945 ;
		RECT	14.565 385.505 14.615 385.635 ;
		RECT	19.885 385.505 19.935 385.635 ;
		RECT	14.765 385.275 14.815 385.405 ;
		RECT	14.765 387.695 14.815 387.825 ;
		RECT	19.685 385.275 19.735 385.405 ;
		RECT	19.685 387.695 19.735 387.825 ;
		RECT	14.965 385.275 15.015 385.405 ;
		RECT	14.965 387.695 15.015 387.825 ;
		RECT	19.485 385.275 19.535 385.405 ;
		RECT	19.485 387.695 19.535 387.825 ;
		RECT	14.565 388.385 14.615 388.515 ;
		RECT	19.885 388.385 19.935 388.515 ;
		RECT	14.765 388.155 14.815 388.285 ;
		RECT	14.765 390.575 14.815 390.705 ;
		RECT	19.685 388.155 19.735 388.285 ;
		RECT	19.685 390.575 19.735 390.705 ;
		RECT	14.965 388.155 15.015 388.285 ;
		RECT	14.965 390.575 15.015 390.705 ;
		RECT	19.485 388.155 19.535 388.285 ;
		RECT	19.485 390.575 19.535 390.705 ;
		RECT	14.565 391.265 14.615 391.395 ;
		RECT	19.885 391.265 19.935 391.395 ;
		RECT	14.765 391.035 14.815 391.165 ;
		RECT	14.765 393.455 14.815 393.585 ;
		RECT	19.685 391.035 19.735 391.165 ;
		RECT	19.685 393.455 19.735 393.585 ;
		RECT	14.965 391.035 15.015 391.165 ;
		RECT	14.965 393.455 15.015 393.585 ;
		RECT	19.485 391.035 19.535 391.165 ;
		RECT	19.485 393.455 19.535 393.585 ;
		RECT	14.565 394.145 14.615 394.275 ;
		RECT	19.885 394.145 19.935 394.275 ;
		RECT	14.765 393.915 14.815 394.045 ;
		RECT	14.765 396.335 14.815 396.465 ;
		RECT	19.685 393.915 19.735 394.045 ;
		RECT	19.685 396.335 19.735 396.465 ;
		RECT	14.965 393.915 15.015 394.045 ;
		RECT	14.965 396.335 15.015 396.465 ;
		RECT	19.485 393.915 19.535 394.045 ;
		RECT	19.485 396.335 19.535 396.465 ;
		RECT	14.565 397.025 14.615 397.155 ;
		RECT	19.885 397.025 19.935 397.155 ;
		RECT	14.765 396.795 14.815 396.925 ;
		RECT	14.765 399.215 14.815 399.345 ;
		RECT	19.685 396.795 19.735 396.925 ;
		RECT	19.685 399.215 19.735 399.345 ;
		RECT	14.965 396.795 15.015 396.925 ;
		RECT	14.965 399.215 15.015 399.345 ;
		RECT	19.485 396.795 19.535 396.925 ;
		RECT	19.485 399.215 19.535 399.345 ;
		RECT	14.565 399.905 14.615 400.035 ;
		RECT	19.885 399.905 19.935 400.035 ;
		RECT	14.765 399.675 14.815 399.805 ;
		RECT	14.765 402.095 14.815 402.225 ;
		RECT	19.685 399.675 19.735 399.805 ;
		RECT	19.685 402.095 19.735 402.225 ;
		RECT	14.965 399.675 15.015 399.805 ;
		RECT	14.965 402.095 15.015 402.225 ;
		RECT	19.485 399.675 19.535 399.805 ;
		RECT	19.485 402.095 19.535 402.225 ;
		RECT	14.565 247.265 14.615 247.395 ;
		RECT	19.885 247.265 19.935 247.395 ;
		RECT	14.765 247.035 14.815 247.165 ;
		RECT	14.765 249.455 14.815 249.585 ;
		RECT	19.685 247.035 19.735 247.165 ;
		RECT	19.685 249.455 19.735 249.585 ;
		RECT	14.965 247.035 15.015 247.165 ;
		RECT	14.965 249.455 15.015 249.585 ;
		RECT	19.485 247.035 19.535 247.165 ;
		RECT	19.485 249.455 19.535 249.585 ;
		RECT	14.565 402.785 14.615 402.915 ;
		RECT	19.885 402.785 19.935 402.915 ;
		RECT	14.765 402.555 14.815 402.685 ;
		RECT	14.765 404.975 14.815 405.105 ;
		RECT	19.685 402.555 19.735 402.685 ;
		RECT	19.685 404.975 19.735 405.105 ;
		RECT	14.965 402.555 15.015 402.685 ;
		RECT	14.965 404.975 15.015 405.105 ;
		RECT	19.485 402.555 19.535 402.685 ;
		RECT	19.485 404.975 19.535 405.105 ;
		RECT	14.565 405.665 14.615 405.795 ;
		RECT	19.885 405.665 19.935 405.795 ;
		RECT	14.765 405.435 14.815 405.565 ;
		RECT	14.765 407.855 14.815 407.985 ;
		RECT	19.685 405.435 19.735 405.565 ;
		RECT	19.685 407.855 19.735 407.985 ;
		RECT	14.965 405.435 15.015 405.565 ;
		RECT	14.965 407.855 15.015 407.985 ;
		RECT	19.485 405.435 19.535 405.565 ;
		RECT	19.485 407.855 19.535 407.985 ;
		RECT	14.565 408.545 14.615 408.675 ;
		RECT	19.885 408.545 19.935 408.675 ;
		RECT	14.765 408.315 14.815 408.445 ;
		RECT	14.765 410.735 14.815 410.865 ;
		RECT	19.685 408.315 19.735 408.445 ;
		RECT	19.685 410.735 19.735 410.865 ;
		RECT	14.965 408.315 15.015 408.445 ;
		RECT	14.965 410.735 15.015 410.865 ;
		RECT	19.485 408.315 19.535 408.445 ;
		RECT	19.485 410.735 19.535 410.865 ;
		RECT	14.565 250.145 14.615 250.275 ;
		RECT	19.885 250.145 19.935 250.275 ;
		RECT	14.765 249.915 14.815 250.045 ;
		RECT	14.765 252.335 14.815 252.465 ;
		RECT	19.685 249.915 19.735 250.045 ;
		RECT	19.685 252.335 19.735 252.465 ;
		RECT	14.965 249.915 15.015 250.045 ;
		RECT	14.965 252.335 15.015 252.465 ;
		RECT	19.485 249.915 19.535 250.045 ;
		RECT	19.485 252.335 19.535 252.465 ;
		RECT	14.565 253.025 14.615 253.155 ;
		RECT	19.885 253.025 19.935 253.155 ;
		RECT	14.765 252.795 14.815 252.925 ;
		RECT	14.765 255.215 14.815 255.345 ;
		RECT	19.685 252.795 19.735 252.925 ;
		RECT	19.685 255.215 19.735 255.345 ;
		RECT	14.965 252.795 15.015 252.925 ;
		RECT	14.965 255.215 15.015 255.345 ;
		RECT	19.485 252.795 19.535 252.925 ;
		RECT	19.485 255.215 19.535 255.345 ;
		RECT	14.565 255.905 14.615 256.035 ;
		RECT	19.885 255.905 19.935 256.035 ;
		RECT	14.765 255.675 14.815 255.805 ;
		RECT	14.765 258.095 14.815 258.225 ;
		RECT	19.685 255.675 19.735 255.805 ;
		RECT	19.685 258.095 19.735 258.225 ;
		RECT	14.965 255.675 15.015 255.805 ;
		RECT	14.965 258.095 15.015 258.225 ;
		RECT	19.485 255.675 19.535 255.805 ;
		RECT	19.485 258.095 19.535 258.225 ;
		RECT	20.085 232.635 20.265 232.765 ;
		RECT	20.875 232.865 21.055 232.995 ;
		RECT	20.085 235.055 20.265 235.185 ;
		RECT	20.43 235.285 20.48 235.415 ;
		RECT	20.085 258.555 20.265 258.685 ;
		RECT	20.875 258.785 21.055 258.915 ;
		RECT	20.085 260.975 20.265 261.105 ;
		RECT	20.43 261.205 20.48 261.335 ;
		RECT	20.085 261.435 20.265 261.565 ;
		RECT	20.875 261.665 21.055 261.795 ;
		RECT	20.085 263.855 20.265 263.985 ;
		RECT	20.43 264.085 20.48 264.215 ;
		RECT	20.085 264.315 20.265 264.445 ;
		RECT	20.875 264.545 21.055 264.675 ;
		RECT	20.085 266.735 20.265 266.865 ;
		RECT	20.43 266.965 20.48 267.095 ;
		RECT	20.085 267.195 20.265 267.325 ;
		RECT	20.875 267.425 21.055 267.555 ;
		RECT	20.085 269.615 20.265 269.745 ;
		RECT	20.43 269.845 20.48 269.975 ;
		RECT	20.085 270.075 20.265 270.205 ;
		RECT	20.875 270.305 21.055 270.435 ;
		RECT	20.085 272.495 20.265 272.625 ;
		RECT	20.43 272.725 20.48 272.855 ;
		RECT	20.085 272.955 20.265 273.085 ;
		RECT	20.875 273.185 21.055 273.315 ;
		RECT	20.085 275.375 20.265 275.505 ;
		RECT	20.43 275.605 20.48 275.735 ;
		RECT	20.085 275.835 20.265 275.965 ;
		RECT	20.875 276.065 21.055 276.195 ;
		RECT	20.085 278.255 20.265 278.385 ;
		RECT	20.43 278.485 20.48 278.615 ;
		RECT	20.085 278.715 20.265 278.845 ;
		RECT	20.875 278.945 21.055 279.075 ;
		RECT	20.085 281.135 20.265 281.265 ;
		RECT	20.43 281.365 20.48 281.495 ;
		RECT	20.085 281.595 20.265 281.725 ;
		RECT	20.875 281.825 21.055 281.955 ;
		RECT	20.085 284.015 20.265 284.145 ;
		RECT	20.43 284.245 20.48 284.375 ;
		RECT	20.085 284.475 20.265 284.605 ;
		RECT	20.875 284.705 21.055 284.835 ;
		RECT	20.085 286.895 20.265 287.025 ;
		RECT	20.43 287.125 20.48 287.255 ;
		RECT	20.085 235.515 20.265 235.645 ;
		RECT	20.875 235.745 21.055 235.875 ;
		RECT	20.085 237.935 20.265 238.065 ;
		RECT	20.43 238.165 20.48 238.295 ;
		RECT	20.085 287.355 20.265 287.485 ;
		RECT	20.875 287.585 21.055 287.715 ;
		RECT	20.085 289.775 20.265 289.905 ;
		RECT	20.43 290.005 20.48 290.135 ;
		RECT	20.085 290.235 20.265 290.365 ;
		RECT	20.875 290.465 21.055 290.595 ;
		RECT	20.085 292.655 20.265 292.785 ;
		RECT	20.43 292.885 20.48 293.015 ;
		RECT	20.085 293.115 20.265 293.245 ;
		RECT	20.875 293.345 21.055 293.475 ;
		RECT	20.085 295.535 20.265 295.665 ;
		RECT	20.43 295.765 20.48 295.895 ;
		RECT	20.085 295.995 20.265 296.125 ;
		RECT	20.875 296.225 21.055 296.355 ;
		RECT	20.085 298.415 20.265 298.545 ;
		RECT	20.43 298.645 20.48 298.775 ;
		RECT	20.085 298.875 20.265 299.005 ;
		RECT	20.875 299.105 21.055 299.235 ;
		RECT	20.085 301.295 20.265 301.425 ;
		RECT	20.43 301.525 20.48 301.655 ;
		RECT	20.085 301.755 20.265 301.885 ;
		RECT	20.875 301.985 21.055 302.115 ;
		RECT	20.085 304.175 20.265 304.305 ;
		RECT	20.43 304.405 20.48 304.535 ;
		RECT	20.085 304.635 20.265 304.765 ;
		RECT	20.875 304.865 21.055 304.995 ;
		RECT	20.085 307.055 20.265 307.185 ;
		RECT	20.43 307.285 20.48 307.415 ;
		RECT	20.085 307.515 20.265 307.645 ;
		RECT	20.875 307.745 21.055 307.875 ;
		RECT	20.085 309.935 20.265 310.065 ;
		RECT	20.43 310.165 20.48 310.295 ;
		RECT	20.085 310.395 20.265 310.525 ;
		RECT	20.875 310.625 21.055 310.755 ;
		RECT	20.085 312.815 20.265 312.945 ;
		RECT	20.43 313.045 20.48 313.175 ;
		RECT	20.085 313.275 20.265 313.405 ;
		RECT	20.875 313.505 21.055 313.635 ;
		RECT	20.085 315.695 20.265 315.825 ;
		RECT	20.43 315.925 20.48 316.055 ;
		RECT	20.085 238.395 20.265 238.525 ;
		RECT	20.875 238.625 21.055 238.755 ;
		RECT	20.085 240.815 20.265 240.945 ;
		RECT	20.43 241.045 20.48 241.175 ;
		RECT	20.085 316.155 20.265 316.285 ;
		RECT	20.875 316.385 21.055 316.515 ;
		RECT	20.085 318.575 20.265 318.705 ;
		RECT	20.43 318.805 20.48 318.935 ;
		RECT	20.085 319.035 20.265 319.165 ;
		RECT	20.875 319.265 21.055 319.395 ;
		RECT	20.085 321.455 20.265 321.585 ;
		RECT	20.43 321.685 20.48 321.815 ;
		RECT	20.085 321.915 20.265 322.045 ;
		RECT	20.875 322.145 21.055 322.275 ;
		RECT	20.085 324.335 20.265 324.465 ;
		RECT	20.43 324.565 20.48 324.695 ;
		RECT	20.085 324.795 20.265 324.925 ;
		RECT	20.875 325.025 21.055 325.155 ;
		RECT	20.085 327.215 20.265 327.345 ;
		RECT	20.43 327.445 20.48 327.575 ;
		RECT	20.085 327.675 20.265 327.805 ;
		RECT	20.875 327.905 21.055 328.035 ;
		RECT	20.085 330.095 20.265 330.225 ;
		RECT	20.43 330.325 20.48 330.455 ;
		RECT	20.085 330.555 20.265 330.685 ;
		RECT	20.875 330.785 21.055 330.915 ;
		RECT	20.085 332.975 20.265 333.105 ;
		RECT	20.43 333.205 20.48 333.335 ;
		RECT	20.085 333.435 20.265 333.565 ;
		RECT	20.875 333.665 21.055 333.795 ;
		RECT	20.085 335.855 20.265 335.985 ;
		RECT	20.43 336.085 20.48 336.215 ;
		RECT	20.085 336.315 20.265 336.445 ;
		RECT	20.875 336.545 21.055 336.675 ;
		RECT	20.085 338.735 20.265 338.865 ;
		RECT	20.43 338.965 20.48 339.095 ;
		RECT	20.085 339.195 20.265 339.325 ;
		RECT	20.875 339.425 21.055 339.555 ;
		RECT	20.085 341.615 20.265 341.745 ;
		RECT	20.43 341.845 20.48 341.975 ;
		RECT	20.085 342.075 20.265 342.205 ;
		RECT	20.875 342.305 21.055 342.435 ;
		RECT	20.085 344.495 20.265 344.625 ;
		RECT	20.43 344.725 20.48 344.855 ;
		RECT	20.085 241.275 20.265 241.405 ;
		RECT	20.875 241.505 21.055 241.635 ;
		RECT	20.085 243.695 20.265 243.825 ;
		RECT	20.43 243.925 20.48 244.055 ;
		RECT	20.085 344.955 20.265 345.085 ;
		RECT	20.875 345.185 21.055 345.315 ;
		RECT	20.085 347.375 20.265 347.505 ;
		RECT	20.43 347.605 20.48 347.735 ;
		RECT	20.085 347.835 20.265 347.965 ;
		RECT	20.875 348.065 21.055 348.195 ;
		RECT	20.085 350.255 20.265 350.385 ;
		RECT	20.43 350.485 20.48 350.615 ;
		RECT	20.085 350.715 20.265 350.845 ;
		RECT	20.875 350.945 21.055 351.075 ;
		RECT	20.085 353.135 20.265 353.265 ;
		RECT	20.43 353.365 20.48 353.495 ;
		RECT	20.085 353.595 20.265 353.725 ;
		RECT	20.875 353.825 21.055 353.955 ;
		RECT	20.085 356.015 20.265 356.145 ;
		RECT	20.43 356.245 20.48 356.375 ;
		RECT	20.085 356.475 20.265 356.605 ;
		RECT	20.875 356.705 21.055 356.835 ;
		RECT	20.085 358.895 20.265 359.025 ;
		RECT	20.43 359.125 20.48 359.255 ;
		RECT	20.085 359.355 20.265 359.485 ;
		RECT	20.875 359.585 21.055 359.715 ;
		RECT	20.085 361.775 20.265 361.905 ;
		RECT	20.43 362.005 20.48 362.135 ;
		RECT	20.085 362.235 20.265 362.365 ;
		RECT	20.875 362.465 21.055 362.595 ;
		RECT	20.085 364.655 20.265 364.785 ;
		RECT	20.43 364.885 20.48 365.015 ;
		RECT	20.085 365.115 20.265 365.245 ;
		RECT	20.875 365.345 21.055 365.475 ;
		RECT	20.085 367.535 20.265 367.665 ;
		RECT	20.43 367.765 20.48 367.895 ;
		RECT	20.085 367.995 20.265 368.125 ;
		RECT	20.875 368.225 21.055 368.355 ;
		RECT	20.085 370.415 20.265 370.545 ;
		RECT	20.43 370.645 20.48 370.775 ;
		RECT	20.085 370.875 20.265 371.005 ;
		RECT	20.875 371.105 21.055 371.235 ;
		RECT	20.085 373.295 20.265 373.425 ;
		RECT	20.43 373.525 20.48 373.655 ;
		RECT	20.085 244.155 20.265 244.285 ;
		RECT	20.875 244.385 21.055 244.515 ;
		RECT	20.085 246.575 20.265 246.705 ;
		RECT	20.43 246.805 20.48 246.935 ;
		RECT	20.085 373.755 20.265 373.885 ;
		RECT	20.875 373.985 21.055 374.115 ;
		RECT	20.085 376.175 20.265 376.305 ;
		RECT	20.43 376.405 20.48 376.535 ;
		RECT	20.085 376.635 20.265 376.765 ;
		RECT	20.875 376.865 21.055 376.995 ;
		RECT	20.085 379.055 20.265 379.185 ;
		RECT	20.43 379.285 20.48 379.415 ;
		RECT	20.085 379.515 20.265 379.645 ;
		RECT	20.875 379.745 21.055 379.875 ;
		RECT	20.085 381.935 20.265 382.065 ;
		RECT	20.43 382.165 20.48 382.295 ;
		RECT	20.085 382.395 20.265 382.525 ;
		RECT	20.875 382.625 21.055 382.755 ;
		RECT	20.085 384.815 20.265 384.945 ;
		RECT	20.43 385.045 20.48 385.175 ;
		RECT	20.085 385.275 20.265 385.405 ;
		RECT	20.875 385.505 21.055 385.635 ;
		RECT	20.085 387.695 20.265 387.825 ;
		RECT	20.43 387.925 20.48 388.055 ;
		RECT	20.085 388.155 20.265 388.285 ;
		RECT	20.875 388.385 21.055 388.515 ;
		RECT	20.085 390.575 20.265 390.705 ;
		RECT	20.43 390.805 20.48 390.935 ;
		RECT	20.085 391.035 20.265 391.165 ;
		RECT	20.875 391.265 21.055 391.395 ;
		RECT	20.085 393.455 20.265 393.585 ;
		RECT	20.43 393.685 20.48 393.815 ;
		RECT	20.085 393.915 20.265 394.045 ;
		RECT	20.875 394.145 21.055 394.275 ;
		RECT	20.085 396.335 20.265 396.465 ;
		RECT	20.43 396.565 20.48 396.695 ;
		RECT	20.085 396.795 20.265 396.925 ;
		RECT	20.875 397.025 21.055 397.155 ;
		RECT	20.085 399.215 20.265 399.345 ;
		RECT	20.43 399.445 20.48 399.575 ;
		RECT	20.085 399.675 20.265 399.805 ;
		RECT	20.875 399.905 21.055 400.035 ;
		RECT	20.085 402.095 20.265 402.225 ;
		RECT	20.43 402.325 20.48 402.455 ;
		RECT	20.085 247.035 20.265 247.165 ;
		RECT	20.875 247.265 21.055 247.395 ;
		RECT	20.085 249.455 20.265 249.585 ;
		RECT	20.43 249.685 20.48 249.815 ;
		RECT	20.085 402.555 20.265 402.685 ;
		RECT	20.875 402.785 21.055 402.915 ;
		RECT	20.085 404.975 20.265 405.105 ;
		RECT	20.43 405.205 20.48 405.335 ;
		RECT	20.085 405.435 20.265 405.565 ;
		RECT	20.875 405.665 21.055 405.795 ;
		RECT	20.085 407.855 20.265 407.985 ;
		RECT	20.43 408.085 20.48 408.215 ;
		RECT	20.085 408.315 20.265 408.445 ;
		RECT	20.875 408.545 21.055 408.675 ;
		RECT	20.085 410.735 20.265 410.865 ;
		RECT	20.43 410.965 20.48 411.095 ;
		RECT	20.085 249.915 20.265 250.045 ;
		RECT	20.875 250.145 21.055 250.275 ;
		RECT	20.085 252.335 20.265 252.465 ;
		RECT	20.43 252.565 20.48 252.695 ;
		RECT	20.085 252.795 20.265 252.925 ;
		RECT	20.875 253.025 21.055 253.155 ;
		RECT	20.085 255.215 20.265 255.345 ;
		RECT	20.43 255.445 20.48 255.575 ;
		RECT	20.085 255.675 20.265 255.805 ;
		RECT	20.875 255.905 21.055 256.035 ;
		RECT	20.085 258.095 20.265 258.225 ;
		RECT	20.43 258.325 20.48 258.455 ;
		RECT	20.085 411.195 20.265 411.325 ;
		RECT	20.875 411.425 21.055 411.555 ;
		RECT	20.085 413.615 20.265 413.745 ;
		RECT	20.43 413.845 20.48 413.975 ;
		RECT	20.085 229.755 20.265 229.885 ;
		RECT	20.875 229.985 21.055 230.115 ;
		RECT	20.085 232.175 20.265 232.305 ;
		RECT	20.43 232.405 20.48 232.535 ;
		RECT	6.225 124.955 6.275 125.085 ;
		RECT	7.5 124.955 7.55 125.085 ;
		RECT	9.04 124.955 9.09 125.085 ;
		RECT	9.315 124.955 9.365 125.085 ;
		RECT	11.025 124.955 11.075 125.085 ;
		RECT	12.79 124.955 12.84 125.085 ;
		RECT	7.18 124.725 7.23 124.855 ;
		RECT	14.14 124.725 14.19 124.855 ;
		RECT	8.56 127.375 8.61 127.505 ;
		RECT	10.27 127.375 10.32 127.505 ;
		RECT	8.56 124.955 8.61 125.085 ;
		RECT	10.27 124.955 10.32 125.085 ;
		RECT	6.22 124.495 6.27 124.625 ;
		RECT	7.5 124.495 7.55 124.625 ;
		RECT	9.04 124.495 9.09 124.625 ;
		RECT	9.315 124.495 9.365 124.625 ;
		RECT	9.72 124.495 9.77 124.625 ;
		RECT	11.025 124.495 11.075 124.625 ;
		RECT	12.79 124.495 12.84 124.625 ;
		RECT	6.225 122.075 6.275 122.205 ;
		RECT	7.5 122.075 7.55 122.205 ;
		RECT	9.04 122.075 9.09 122.205 ;
		RECT	9.315 122.075 9.365 122.205 ;
		RECT	11.025 122.075 11.075 122.205 ;
		RECT	12.79 122.075 12.84 122.205 ;
		RECT	7.18 121.845 7.23 121.975 ;
		RECT	14.14 121.845 14.19 121.975 ;
		RECT	8.56 124.495 8.61 124.625 ;
		RECT	10.27 124.495 10.32 124.625 ;
		RECT	8.56 122.075 8.61 122.205 ;
		RECT	10.27 122.075 10.32 122.205 ;
		RECT	6.22 121.615 6.27 121.745 ;
		RECT	7.5 121.615 7.55 121.745 ;
		RECT	9.04 121.615 9.09 121.745 ;
		RECT	9.315 121.615 9.365 121.745 ;
		RECT	9.72 121.615 9.77 121.745 ;
		RECT	11.025 121.615 11.075 121.745 ;
		RECT	12.79 121.615 12.84 121.745 ;
		RECT	6.225 119.195 6.275 119.325 ;
		RECT	7.5 119.195 7.55 119.325 ;
		RECT	9.04 119.195 9.09 119.325 ;
		RECT	9.315 119.195 9.365 119.325 ;
		RECT	11.025 119.195 11.075 119.325 ;
		RECT	12.79 119.195 12.84 119.325 ;
		RECT	7.18 118.965 7.23 119.095 ;
		RECT	14.14 118.965 14.19 119.095 ;
		RECT	8.56 121.615 8.61 121.745 ;
		RECT	10.27 121.615 10.32 121.745 ;
		RECT	8.56 119.195 8.61 119.325 ;
		RECT	10.27 119.195 10.32 119.325 ;
		RECT	6.22 118.735 6.27 118.865 ;
		RECT	7.5 118.735 7.55 118.865 ;
		RECT	9.04 118.735 9.09 118.865 ;
		RECT	9.315 118.735 9.365 118.865 ;
		RECT	9.72 118.735 9.77 118.865 ;
		RECT	11.025 118.735 11.075 118.865 ;
		RECT	12.79 118.735 12.84 118.865 ;
		RECT	6.225 116.315 6.275 116.445 ;
		RECT	7.5 116.315 7.55 116.445 ;
		RECT	9.04 116.315 9.09 116.445 ;
		RECT	9.315 116.315 9.365 116.445 ;
		RECT	11.025 116.315 11.075 116.445 ;
		RECT	12.79 116.315 12.84 116.445 ;
		RECT	7.18 116.085 7.23 116.215 ;
		RECT	14.14 116.085 14.19 116.215 ;
		RECT	8.56 118.735 8.61 118.865 ;
		RECT	10.27 118.735 10.32 118.865 ;
		RECT	8.56 116.315 8.61 116.445 ;
		RECT	10.27 116.315 10.32 116.445 ;
		RECT	6.22 115.855 6.27 115.985 ;
		RECT	7.5 115.855 7.55 115.985 ;
		RECT	9.04 115.855 9.09 115.985 ;
		RECT	9.315 115.855 9.365 115.985 ;
		RECT	9.72 115.855 9.77 115.985 ;
		RECT	11.025 115.855 11.075 115.985 ;
		RECT	12.79 115.855 12.84 115.985 ;
		RECT	6.225 113.435 6.275 113.565 ;
		RECT	7.5 113.435 7.55 113.565 ;
		RECT	9.04 113.435 9.09 113.565 ;
		RECT	9.315 113.435 9.365 113.565 ;
		RECT	11.025 113.435 11.075 113.565 ;
		RECT	12.79 113.435 12.84 113.565 ;
		RECT	7.18 113.205 7.23 113.335 ;
		RECT	14.14 113.205 14.19 113.335 ;
		RECT	8.56 115.855 8.61 115.985 ;
		RECT	10.27 115.855 10.32 115.985 ;
		RECT	8.56 113.435 8.61 113.565 ;
		RECT	10.27 113.435 10.32 113.565 ;
		RECT	6.22 112.975 6.27 113.105 ;
		RECT	7.5 112.975 7.55 113.105 ;
		RECT	9.04 112.975 9.09 113.105 ;
		RECT	9.315 112.975 9.365 113.105 ;
		RECT	9.72 112.975 9.77 113.105 ;
		RECT	11.025 112.975 11.075 113.105 ;
		RECT	12.79 112.975 12.84 113.105 ;
		RECT	6.225 110.555 6.275 110.685 ;
		RECT	7.5 110.555 7.55 110.685 ;
		RECT	9.04 110.555 9.09 110.685 ;
		RECT	9.315 110.555 9.365 110.685 ;
		RECT	11.025 110.555 11.075 110.685 ;
		RECT	12.79 110.555 12.84 110.685 ;
		RECT	7.18 110.325 7.23 110.455 ;
		RECT	14.14 110.325 14.19 110.455 ;
		RECT	8.56 112.975 8.61 113.105 ;
		RECT	10.27 112.975 10.32 113.105 ;
		RECT	8.56 110.555 8.61 110.685 ;
		RECT	10.27 110.555 10.32 110.685 ;
		RECT	6.22 110.095 6.27 110.225 ;
		RECT	7.5 110.095 7.55 110.225 ;
		RECT	9.04 110.095 9.09 110.225 ;
		RECT	9.315 110.095 9.365 110.225 ;
		RECT	9.72 110.095 9.77 110.225 ;
		RECT	11.025 110.095 11.075 110.225 ;
		RECT	12.79 110.095 12.84 110.225 ;
		RECT	6.225 107.675 6.275 107.805 ;
		RECT	7.5 107.675 7.55 107.805 ;
		RECT	9.04 107.675 9.09 107.805 ;
		RECT	9.315 107.675 9.365 107.805 ;
		RECT	11.025 107.675 11.075 107.805 ;
		RECT	12.79 107.675 12.84 107.805 ;
		RECT	7.18 107.445 7.23 107.575 ;
		RECT	14.14 107.445 14.19 107.575 ;
		RECT	8.56 110.095 8.61 110.225 ;
		RECT	10.27 110.095 10.32 110.225 ;
		RECT	8.56 107.675 8.61 107.805 ;
		RECT	10.27 107.675 10.32 107.805 ;
		RECT	6.22 107.215 6.27 107.345 ;
		RECT	7.5 107.215 7.55 107.345 ;
		RECT	9.04 107.215 9.09 107.345 ;
		RECT	9.315 107.215 9.365 107.345 ;
		RECT	9.72 107.215 9.77 107.345 ;
		RECT	11.025 107.215 11.075 107.345 ;
		RECT	12.79 107.215 12.84 107.345 ;
		RECT	6.225 104.795 6.275 104.925 ;
		RECT	7.5 104.795 7.55 104.925 ;
		RECT	9.04 104.795 9.09 104.925 ;
		RECT	9.315 104.795 9.365 104.925 ;
		RECT	11.025 104.795 11.075 104.925 ;
		RECT	12.79 104.795 12.84 104.925 ;
		RECT	7.18 104.565 7.23 104.695 ;
		RECT	14.14 104.565 14.19 104.695 ;
		RECT	8.56 107.215 8.61 107.345 ;
		RECT	10.27 107.215 10.32 107.345 ;
		RECT	8.56 104.795 8.61 104.925 ;
		RECT	10.27 104.795 10.32 104.925 ;
		RECT	6.22 104.335 6.27 104.465 ;
		RECT	7.5 104.335 7.55 104.465 ;
		RECT	9.04 104.335 9.09 104.465 ;
		RECT	9.315 104.335 9.365 104.465 ;
		RECT	9.72 104.335 9.77 104.465 ;
		RECT	11.025 104.335 11.075 104.465 ;
		RECT	12.79 104.335 12.84 104.465 ;
		RECT	6.225 101.915 6.275 102.045 ;
		RECT	7.5 101.915 7.55 102.045 ;
		RECT	9.04 101.915 9.09 102.045 ;
		RECT	9.315 101.915 9.365 102.045 ;
		RECT	11.025 101.915 11.075 102.045 ;
		RECT	12.79 101.915 12.84 102.045 ;
		RECT	7.18 101.685 7.23 101.815 ;
		RECT	14.14 101.685 14.19 101.815 ;
		RECT	8.56 104.335 8.61 104.465 ;
		RECT	10.27 104.335 10.32 104.465 ;
		RECT	8.56 101.915 8.61 102.045 ;
		RECT	10.27 101.915 10.32 102.045 ;
		RECT	6.22 101.455 6.27 101.585 ;
		RECT	7.5 101.455 7.55 101.585 ;
		RECT	9.04 101.455 9.09 101.585 ;
		RECT	9.315 101.455 9.365 101.585 ;
		RECT	9.72 101.455 9.77 101.585 ;
		RECT	11.025 101.455 11.075 101.585 ;
		RECT	12.79 101.455 12.84 101.585 ;
		RECT	6.225 99.035 6.275 99.165 ;
		RECT	7.5 99.035 7.55 99.165 ;
		RECT	9.04 99.035 9.09 99.165 ;
		RECT	9.315 99.035 9.365 99.165 ;
		RECT	11.025 99.035 11.075 99.165 ;
		RECT	12.79 99.035 12.84 99.165 ;
		RECT	7.18 98.805 7.23 98.935 ;
		RECT	14.14 98.805 14.19 98.935 ;
		RECT	8.56 101.455 8.61 101.585 ;
		RECT	10.27 101.455 10.32 101.585 ;
		RECT	8.56 99.035 8.61 99.165 ;
		RECT	10.27 99.035 10.32 99.165 ;
		RECT	6.22 98.575 6.27 98.705 ;
		RECT	7.5 98.575 7.55 98.705 ;
		RECT	9.04 98.575 9.09 98.705 ;
		RECT	9.315 98.575 9.365 98.705 ;
		RECT	9.72 98.575 9.77 98.705 ;
		RECT	11.025 98.575 11.075 98.705 ;
		RECT	12.79 98.575 12.84 98.705 ;
		RECT	6.225 96.155 6.275 96.285 ;
		RECT	7.5 96.155 7.55 96.285 ;
		RECT	9.04 96.155 9.09 96.285 ;
		RECT	9.315 96.155 9.365 96.285 ;
		RECT	11.025 96.155 11.075 96.285 ;
		RECT	12.79 96.155 12.84 96.285 ;
		RECT	7.18 95.925 7.23 96.055 ;
		RECT	14.14 95.925 14.19 96.055 ;
		RECT	8.56 98.575 8.61 98.705 ;
		RECT	10.27 98.575 10.32 98.705 ;
		RECT	8.56 96.155 8.61 96.285 ;
		RECT	10.27 96.155 10.32 96.285 ;
		RECT	6.22 95.695 6.27 95.825 ;
		RECT	7.5 95.695 7.55 95.825 ;
		RECT	9.04 95.695 9.09 95.825 ;
		RECT	9.315 95.695 9.365 95.825 ;
		RECT	9.72 95.695 9.77 95.825 ;
		RECT	11.025 95.695 11.075 95.825 ;
		RECT	12.79 95.695 12.84 95.825 ;
		RECT	6.225 93.275 6.275 93.405 ;
		RECT	7.5 93.275 7.55 93.405 ;
		RECT	9.04 93.275 9.09 93.405 ;
		RECT	9.315 93.275 9.365 93.405 ;
		RECT	11.025 93.275 11.075 93.405 ;
		RECT	12.79 93.275 12.84 93.405 ;
		RECT	7.18 93.045 7.23 93.175 ;
		RECT	14.14 93.045 14.19 93.175 ;
		RECT	8.56 95.695 8.61 95.825 ;
		RECT	10.27 95.695 10.32 95.825 ;
		RECT	8.56 93.275 8.61 93.405 ;
		RECT	10.27 93.275 10.32 93.405 ;
		RECT	6.22 92.815 6.27 92.945 ;
		RECT	7.5 92.815 7.55 92.945 ;
		RECT	9.04 92.815 9.09 92.945 ;
		RECT	9.315 92.815 9.365 92.945 ;
		RECT	9.72 92.815 9.77 92.945 ;
		RECT	11.025 92.815 11.075 92.945 ;
		RECT	12.79 92.815 12.84 92.945 ;
		RECT	6.225 90.395 6.275 90.525 ;
		RECT	7.5 90.395 7.55 90.525 ;
		RECT	9.04 90.395 9.09 90.525 ;
		RECT	9.315 90.395 9.365 90.525 ;
		RECT	11.025 90.395 11.075 90.525 ;
		RECT	12.79 90.395 12.84 90.525 ;
		RECT	7.18 90.165 7.23 90.295 ;
		RECT	14.14 90.165 14.19 90.295 ;
		RECT	8.56 92.815 8.61 92.945 ;
		RECT	10.27 92.815 10.32 92.945 ;
		RECT	8.56 90.395 8.61 90.525 ;
		RECT	10.27 90.395 10.32 90.525 ;
		RECT	6.22 89.935 6.27 90.065 ;
		RECT	7.5 89.935 7.55 90.065 ;
		RECT	9.04 89.935 9.09 90.065 ;
		RECT	9.315 89.935 9.365 90.065 ;
		RECT	9.72 89.935 9.77 90.065 ;
		RECT	11.025 89.935 11.075 90.065 ;
		RECT	12.79 89.935 12.84 90.065 ;
		RECT	6.225 87.515 6.275 87.645 ;
		RECT	7.5 87.515 7.55 87.645 ;
		RECT	9.04 87.515 9.09 87.645 ;
		RECT	9.315 87.515 9.365 87.645 ;
		RECT	11.025 87.515 11.075 87.645 ;
		RECT	12.79 87.515 12.84 87.645 ;
		RECT	7.18 87.285 7.23 87.415 ;
		RECT	14.14 87.285 14.19 87.415 ;
		RECT	8.56 89.935 8.61 90.065 ;
		RECT	10.27 89.935 10.32 90.065 ;
		RECT	8.56 87.515 8.61 87.645 ;
		RECT	10.27 87.515 10.32 87.645 ;
		RECT	6.22 87.055 6.27 87.185 ;
		RECT	7.5 87.055 7.55 87.185 ;
		RECT	9.04 87.055 9.09 87.185 ;
		RECT	9.315 87.055 9.365 87.185 ;
		RECT	9.72 87.055 9.77 87.185 ;
		RECT	11.025 87.055 11.075 87.185 ;
		RECT	12.79 87.055 12.84 87.185 ;
		RECT	6.225 84.635 6.275 84.765 ;
		RECT	7.5 84.635 7.55 84.765 ;
		RECT	9.04 84.635 9.09 84.765 ;
		RECT	9.315 84.635 9.365 84.765 ;
		RECT	11.025 84.635 11.075 84.765 ;
		RECT	12.79 84.635 12.84 84.765 ;
		RECT	7.18 84.405 7.23 84.535 ;
		RECT	14.14 84.405 14.19 84.535 ;
		RECT	8.56 87.055 8.61 87.185 ;
		RECT	10.27 87.055 10.32 87.185 ;
		RECT	8.56 84.635 8.61 84.765 ;
		RECT	10.27 84.635 10.32 84.765 ;
		RECT	6.22 84.175 6.27 84.305 ;
		RECT	7.5 84.175 7.55 84.305 ;
		RECT	9.04 84.175 9.09 84.305 ;
		RECT	9.315 84.175 9.365 84.305 ;
		RECT	9.72 84.175 9.77 84.305 ;
		RECT	11.025 84.175 11.075 84.305 ;
		RECT	12.79 84.175 12.84 84.305 ;
		RECT	6.225 81.755 6.275 81.885 ;
		RECT	7.5 81.755 7.55 81.885 ;
		RECT	9.04 81.755 9.09 81.885 ;
		RECT	9.315 81.755 9.365 81.885 ;
		RECT	11.025 81.755 11.075 81.885 ;
		RECT	12.79 81.755 12.84 81.885 ;
		RECT	7.18 81.525 7.23 81.655 ;
		RECT	14.14 81.525 14.19 81.655 ;
		RECT	8.56 84.175 8.61 84.305 ;
		RECT	10.27 84.175 10.32 84.305 ;
		RECT	8.56 81.755 8.61 81.885 ;
		RECT	10.27 81.755 10.32 81.885 ;
		RECT	6.22 81.295 6.27 81.425 ;
		RECT	7.5 81.295 7.55 81.425 ;
		RECT	9.04 81.295 9.09 81.425 ;
		RECT	9.315 81.295 9.365 81.425 ;
		RECT	9.72 81.295 9.77 81.425 ;
		RECT	11.025 81.295 11.075 81.425 ;
		RECT	12.79 81.295 12.84 81.425 ;
		RECT	6.225 78.875 6.275 79.005 ;
		RECT	7.5 78.875 7.55 79.005 ;
		RECT	9.04 78.875 9.09 79.005 ;
		RECT	9.315 78.875 9.365 79.005 ;
		RECT	11.025 78.875 11.075 79.005 ;
		RECT	12.79 78.875 12.84 79.005 ;
		RECT	7.18 78.645 7.23 78.775 ;
		RECT	14.14 78.645 14.19 78.775 ;
		RECT	8.56 81.295 8.61 81.425 ;
		RECT	10.27 81.295 10.32 81.425 ;
		RECT	8.56 78.875 8.61 79.005 ;
		RECT	10.27 78.875 10.32 79.005 ;
		RECT	6.22 78.415 6.27 78.545 ;
		RECT	7.5 78.415 7.55 78.545 ;
		RECT	9.04 78.415 9.09 78.545 ;
		RECT	9.315 78.415 9.365 78.545 ;
		RECT	9.72 78.415 9.77 78.545 ;
		RECT	11.025 78.415 11.075 78.545 ;
		RECT	12.79 78.415 12.84 78.545 ;
		RECT	6.225 75.995 6.275 76.125 ;
		RECT	7.5 75.995 7.55 76.125 ;
		RECT	9.04 75.995 9.09 76.125 ;
		RECT	9.315 75.995 9.365 76.125 ;
		RECT	11.025 75.995 11.075 76.125 ;
		RECT	12.79 75.995 12.84 76.125 ;
		RECT	7.18 75.765 7.23 75.895 ;
		RECT	14.14 75.765 14.19 75.895 ;
		RECT	8.56 78.415 8.61 78.545 ;
		RECT	10.27 78.415 10.32 78.545 ;
		RECT	8.56 75.995 8.61 76.125 ;
		RECT	10.27 75.995 10.32 76.125 ;
		RECT	6.22 75.535 6.27 75.665 ;
		RECT	7.5 75.535 7.55 75.665 ;
		RECT	9.04 75.535 9.09 75.665 ;
		RECT	9.315 75.535 9.365 75.665 ;
		RECT	9.72 75.535 9.77 75.665 ;
		RECT	11.025 75.535 11.075 75.665 ;
		RECT	12.79 75.535 12.84 75.665 ;
		RECT	6.225 73.115 6.275 73.245 ;
		RECT	7.5 73.115 7.55 73.245 ;
		RECT	9.04 73.115 9.09 73.245 ;
		RECT	9.315 73.115 9.365 73.245 ;
		RECT	11.025 73.115 11.075 73.245 ;
		RECT	12.79 73.115 12.84 73.245 ;
		RECT	7.18 72.885 7.23 73.015 ;
		RECT	14.14 72.885 14.19 73.015 ;
		RECT	8.56 75.535 8.61 75.665 ;
		RECT	10.27 75.535 10.32 75.665 ;
		RECT	8.56 73.115 8.61 73.245 ;
		RECT	10.27 73.115 10.32 73.245 ;
		RECT	6.22 72.655 6.27 72.785 ;
		RECT	7.5 72.655 7.55 72.785 ;
		RECT	9.04 72.655 9.09 72.785 ;
		RECT	9.315 72.655 9.365 72.785 ;
		RECT	9.72 72.655 9.77 72.785 ;
		RECT	11.025 72.655 11.075 72.785 ;
		RECT	12.79 72.655 12.84 72.785 ;
		RECT	6.225 70.235 6.275 70.365 ;
		RECT	7.5 70.235 7.55 70.365 ;
		RECT	9.04 70.235 9.09 70.365 ;
		RECT	9.315 70.235 9.365 70.365 ;
		RECT	11.025 70.235 11.075 70.365 ;
		RECT	12.79 70.235 12.84 70.365 ;
		RECT	7.18 70.005 7.23 70.135 ;
		RECT	14.14 70.005 14.19 70.135 ;
		RECT	8.56 72.655 8.61 72.785 ;
		RECT	10.27 72.655 10.32 72.785 ;
		RECT	8.56 70.235 8.61 70.365 ;
		RECT	10.27 70.235 10.32 70.365 ;
		RECT	6.22 69.775 6.27 69.905 ;
		RECT	7.5 69.775 7.55 69.905 ;
		RECT	9.04 69.775 9.09 69.905 ;
		RECT	9.315 69.775 9.365 69.905 ;
		RECT	9.72 69.775 9.77 69.905 ;
		RECT	11.025 69.775 11.075 69.905 ;
		RECT	12.79 69.775 12.84 69.905 ;
		RECT	6.225 67.355 6.275 67.485 ;
		RECT	7.5 67.355 7.55 67.485 ;
		RECT	9.04 67.355 9.09 67.485 ;
		RECT	9.315 67.355 9.365 67.485 ;
		RECT	11.025 67.355 11.075 67.485 ;
		RECT	12.79 67.355 12.84 67.485 ;
		RECT	7.18 67.125 7.23 67.255 ;
		RECT	14.14 67.125 14.19 67.255 ;
		RECT	8.56 69.775 8.61 69.905 ;
		RECT	10.27 69.775 10.32 69.905 ;
		RECT	8.56 67.355 8.61 67.485 ;
		RECT	10.27 67.355 10.32 67.485 ;
		RECT	6.22 66.895 6.27 67.025 ;
		RECT	7.5 66.895 7.55 67.025 ;
		RECT	9.04 66.895 9.09 67.025 ;
		RECT	9.315 66.895 9.365 67.025 ;
		RECT	9.72 66.895 9.77 67.025 ;
		RECT	11.025 66.895 11.075 67.025 ;
		RECT	12.79 66.895 12.84 67.025 ;
		RECT	6.225 64.475 6.275 64.605 ;
		RECT	7.5 64.475 7.55 64.605 ;
		RECT	9.04 64.475 9.09 64.605 ;
		RECT	9.315 64.475 9.365 64.605 ;
		RECT	11.025 64.475 11.075 64.605 ;
		RECT	12.79 64.475 12.84 64.605 ;
		RECT	7.18 64.245 7.23 64.375 ;
		RECT	14.14 64.245 14.19 64.375 ;
		RECT	8.56 66.895 8.61 67.025 ;
		RECT	10.27 66.895 10.32 67.025 ;
		RECT	8.56 64.475 8.61 64.605 ;
		RECT	10.27 64.475 10.32 64.605 ;
		RECT	6.22 64.015 6.27 64.145 ;
		RECT	7.5 64.015 7.55 64.145 ;
		RECT	9.04 64.015 9.09 64.145 ;
		RECT	9.315 64.015 9.365 64.145 ;
		RECT	9.72 64.015 9.77 64.145 ;
		RECT	11.025 64.015 11.075 64.145 ;
		RECT	12.79 64.015 12.84 64.145 ;
		RECT	6.225 61.595 6.275 61.725 ;
		RECT	7.5 61.595 7.55 61.725 ;
		RECT	9.04 61.595 9.09 61.725 ;
		RECT	9.315 61.595 9.365 61.725 ;
		RECT	11.025 61.595 11.075 61.725 ;
		RECT	12.79 61.595 12.84 61.725 ;
		RECT	7.18 61.365 7.23 61.495 ;
		RECT	14.14 61.365 14.19 61.495 ;
		RECT	8.56 64.015 8.61 64.145 ;
		RECT	10.27 64.015 10.32 64.145 ;
		RECT	8.56 61.595 8.61 61.725 ;
		RECT	10.27 61.595 10.32 61.725 ;
		RECT	6.22 61.135 6.27 61.265 ;
		RECT	7.5 61.135 7.55 61.265 ;
		RECT	9.04 61.135 9.09 61.265 ;
		RECT	9.315 61.135 9.365 61.265 ;
		RECT	9.72 61.135 9.77 61.265 ;
		RECT	11.025 61.135 11.075 61.265 ;
		RECT	12.79 61.135 12.84 61.265 ;
		RECT	6.225 58.715 6.275 58.845 ;
		RECT	7.5 58.715 7.55 58.845 ;
		RECT	9.04 58.715 9.09 58.845 ;
		RECT	9.315 58.715 9.365 58.845 ;
		RECT	11.025 58.715 11.075 58.845 ;
		RECT	12.79 58.715 12.84 58.845 ;
		RECT	7.18 58.485 7.23 58.615 ;
		RECT	14.14 58.485 14.19 58.615 ;
		RECT	8.56 61.135 8.61 61.265 ;
		RECT	10.27 61.135 10.32 61.265 ;
		RECT	8.56 58.715 8.61 58.845 ;
		RECT	10.27 58.715 10.32 58.845 ;
		RECT	6.22 58.255 6.27 58.385 ;
		RECT	7.5 58.255 7.55 58.385 ;
		RECT	9.04 58.255 9.09 58.385 ;
		RECT	9.315 58.255 9.365 58.385 ;
		RECT	9.72 58.255 9.77 58.385 ;
		RECT	11.025 58.255 11.075 58.385 ;
		RECT	12.79 58.255 12.84 58.385 ;
		RECT	6.225 55.835 6.275 55.965 ;
		RECT	7.5 55.835 7.55 55.965 ;
		RECT	9.04 55.835 9.09 55.965 ;
		RECT	9.315 55.835 9.365 55.965 ;
		RECT	11.025 55.835 11.075 55.965 ;
		RECT	12.79 55.835 12.84 55.965 ;
		RECT	7.18 55.605 7.23 55.735 ;
		RECT	14.14 55.605 14.19 55.735 ;
		RECT	8.56 58.255 8.61 58.385 ;
		RECT	10.27 58.255 10.32 58.385 ;
		RECT	8.56 55.835 8.61 55.965 ;
		RECT	10.27 55.835 10.32 55.965 ;
		RECT	6.22 55.375 6.27 55.505 ;
		RECT	7.5 55.375 7.55 55.505 ;
		RECT	9.04 55.375 9.09 55.505 ;
		RECT	9.315 55.375 9.365 55.505 ;
		RECT	9.72 55.375 9.77 55.505 ;
		RECT	11.025 55.375 11.075 55.505 ;
		RECT	12.79 55.375 12.84 55.505 ;
		RECT	6.225 52.955 6.275 53.085 ;
		RECT	7.5 52.955 7.55 53.085 ;
		RECT	9.04 52.955 9.09 53.085 ;
		RECT	9.315 52.955 9.365 53.085 ;
		RECT	11.025 52.955 11.075 53.085 ;
		RECT	12.79 52.955 12.84 53.085 ;
		RECT	7.18 52.725 7.23 52.855 ;
		RECT	14.14 52.725 14.19 52.855 ;
		RECT	8.56 55.375 8.61 55.505 ;
		RECT	10.27 55.375 10.32 55.505 ;
		RECT	8.56 52.955 8.61 53.085 ;
		RECT	10.27 52.955 10.32 53.085 ;
		RECT	6.22 52.495 6.27 52.625 ;
		RECT	7.5 52.495 7.55 52.625 ;
		RECT	9.04 52.495 9.09 52.625 ;
		RECT	9.315 52.495 9.365 52.625 ;
		RECT	9.72 52.495 9.77 52.625 ;
		RECT	11.025 52.495 11.075 52.625 ;
		RECT	12.79 52.495 12.84 52.625 ;
		RECT	6.225 50.075 6.275 50.205 ;
		RECT	7.5 50.075 7.55 50.205 ;
		RECT	9.04 50.075 9.09 50.205 ;
		RECT	9.315 50.075 9.365 50.205 ;
		RECT	11.025 50.075 11.075 50.205 ;
		RECT	12.79 50.075 12.84 50.205 ;
		RECT	7.18 49.845 7.23 49.975 ;
		RECT	14.14 49.845 14.19 49.975 ;
		RECT	8.56 52.495 8.61 52.625 ;
		RECT	10.27 52.495 10.32 52.625 ;
		RECT	8.56 50.075 8.61 50.205 ;
		RECT	10.27 50.075 10.32 50.205 ;
		RECT	6.22 49.615 6.27 49.745 ;
		RECT	7.5 49.615 7.55 49.745 ;
		RECT	9.04 49.615 9.09 49.745 ;
		RECT	9.315 49.615 9.365 49.745 ;
		RECT	9.72 49.615 9.77 49.745 ;
		RECT	11.025 49.615 11.075 49.745 ;
		RECT	12.79 49.615 12.84 49.745 ;
		RECT	6.225 47.195 6.275 47.325 ;
		RECT	7.5 47.195 7.55 47.325 ;
		RECT	9.04 47.195 9.09 47.325 ;
		RECT	9.315 47.195 9.365 47.325 ;
		RECT	11.025 47.195 11.075 47.325 ;
		RECT	12.79 47.195 12.84 47.325 ;
		RECT	7.18 46.965 7.23 47.095 ;
		RECT	14.14 46.965 14.19 47.095 ;
		RECT	8.56 49.615 8.61 49.745 ;
		RECT	10.27 49.615 10.32 49.745 ;
		RECT	8.56 47.195 8.61 47.325 ;
		RECT	10.27 47.195 10.32 47.325 ;
		RECT	6.22 46.735 6.27 46.865 ;
		RECT	7.5 46.735 7.55 46.865 ;
		RECT	9.04 46.735 9.09 46.865 ;
		RECT	9.315 46.735 9.365 46.865 ;
		RECT	9.72 46.735 9.77 46.865 ;
		RECT	11.025 46.735 11.075 46.865 ;
		RECT	12.79 46.735 12.84 46.865 ;
		RECT	6.225 44.315 6.275 44.445 ;
		RECT	7.5 44.315 7.55 44.445 ;
		RECT	9.04 44.315 9.09 44.445 ;
		RECT	9.315 44.315 9.365 44.445 ;
		RECT	11.025 44.315 11.075 44.445 ;
		RECT	12.79 44.315 12.84 44.445 ;
		RECT	7.18 44.085 7.23 44.215 ;
		RECT	14.14 44.085 14.19 44.215 ;
		RECT	8.56 46.735 8.61 46.865 ;
		RECT	10.27 46.735 10.32 46.865 ;
		RECT	8.56 44.315 8.61 44.445 ;
		RECT	10.27 44.315 10.32 44.445 ;
		RECT	6.22 43.855 6.27 43.985 ;
		RECT	7.5 43.855 7.55 43.985 ;
		RECT	9.04 43.855 9.09 43.985 ;
		RECT	9.315 43.855 9.365 43.985 ;
		RECT	9.72 43.855 9.77 43.985 ;
		RECT	11.025 43.855 11.075 43.985 ;
		RECT	12.79 43.855 12.84 43.985 ;
		RECT	6.225 41.435 6.275 41.565 ;
		RECT	7.5 41.435 7.55 41.565 ;
		RECT	9.04 41.435 9.09 41.565 ;
		RECT	9.315 41.435 9.365 41.565 ;
		RECT	11.025 41.435 11.075 41.565 ;
		RECT	12.79 41.435 12.84 41.565 ;
		RECT	7.18 41.205 7.23 41.335 ;
		RECT	14.14 41.205 14.19 41.335 ;
		RECT	8.56 43.855 8.61 43.985 ;
		RECT	10.27 43.855 10.32 43.985 ;
		RECT	8.56 41.435 8.61 41.565 ;
		RECT	10.27 41.435 10.32 41.565 ;
		RECT	6.22 40.975 6.27 41.105 ;
		RECT	7.5 40.975 7.55 41.105 ;
		RECT	9.04 40.975 9.09 41.105 ;
		RECT	9.315 40.975 9.365 41.105 ;
		RECT	9.72 40.975 9.77 41.105 ;
		RECT	11.025 40.975 11.075 41.105 ;
		RECT	12.79 40.975 12.84 41.105 ;
		RECT	6.225 38.555 6.275 38.685 ;
		RECT	7.5 38.555 7.55 38.685 ;
		RECT	9.04 38.555 9.09 38.685 ;
		RECT	9.315 38.555 9.365 38.685 ;
		RECT	11.025 38.555 11.075 38.685 ;
		RECT	12.79 38.555 12.84 38.685 ;
		RECT	7.18 38.325 7.23 38.455 ;
		RECT	14.14 38.325 14.19 38.455 ;
		RECT	8.56 40.975 8.61 41.105 ;
		RECT	10.27 40.975 10.32 41.105 ;
		RECT	8.56 38.555 8.61 38.685 ;
		RECT	10.27 38.555 10.32 38.685 ;
		RECT	6.22 38.095 6.27 38.225 ;
		RECT	7.5 38.095 7.55 38.225 ;
		RECT	9.04 38.095 9.09 38.225 ;
		RECT	9.315 38.095 9.365 38.225 ;
		RECT	9.72 38.095 9.77 38.225 ;
		RECT	11.025 38.095 11.075 38.225 ;
		RECT	12.79 38.095 12.84 38.225 ;
		RECT	6.225 35.675 6.275 35.805 ;
		RECT	7.5 35.675 7.55 35.805 ;
		RECT	9.04 35.675 9.09 35.805 ;
		RECT	9.315 35.675 9.365 35.805 ;
		RECT	11.025 35.675 11.075 35.805 ;
		RECT	12.79 35.675 12.84 35.805 ;
		RECT	7.18 35.445 7.23 35.575 ;
		RECT	14.14 35.445 14.19 35.575 ;
		RECT	8.56 38.095 8.61 38.225 ;
		RECT	10.27 38.095 10.32 38.225 ;
		RECT	8.56 35.675 8.61 35.805 ;
		RECT	10.27 35.675 10.32 35.805 ;
		RECT	6.22 35.215 6.27 35.345 ;
		RECT	7.5 35.215 7.55 35.345 ;
		RECT	9.04 35.215 9.09 35.345 ;
		RECT	9.315 35.215 9.365 35.345 ;
		RECT	9.72 35.215 9.77 35.345 ;
		RECT	11.025 35.215 11.075 35.345 ;
		RECT	12.79 35.215 12.84 35.345 ;
		RECT	6.225 32.795 6.275 32.925 ;
		RECT	7.5 32.795 7.55 32.925 ;
		RECT	9.04 32.795 9.09 32.925 ;
		RECT	9.315 32.795 9.365 32.925 ;
		RECT	11.025 32.795 11.075 32.925 ;
		RECT	12.79 32.795 12.84 32.925 ;
		RECT	7.18 32.565 7.23 32.695 ;
		RECT	14.14 32.565 14.19 32.695 ;
		RECT	8.56 35.215 8.61 35.345 ;
		RECT	10.27 35.215 10.32 35.345 ;
		RECT	8.56 32.795 8.61 32.925 ;
		RECT	10.27 32.795 10.32 32.925 ;
		RECT	6.22 32.335 6.27 32.465 ;
		RECT	7.5 32.335 7.55 32.465 ;
		RECT	9.04 32.335 9.09 32.465 ;
		RECT	9.315 32.335 9.365 32.465 ;
		RECT	9.72 32.335 9.77 32.465 ;
		RECT	11.025 32.335 11.075 32.465 ;
		RECT	12.79 32.335 12.84 32.465 ;
		RECT	6.225 29.915 6.275 30.045 ;
		RECT	7.5 29.915 7.55 30.045 ;
		RECT	9.04 29.915 9.09 30.045 ;
		RECT	9.315 29.915 9.365 30.045 ;
		RECT	11.025 29.915 11.075 30.045 ;
		RECT	12.79 29.915 12.84 30.045 ;
		RECT	7.18 29.685 7.23 29.815 ;
		RECT	14.14 29.685 14.19 29.815 ;
		RECT	8.56 32.335 8.61 32.465 ;
		RECT	10.27 32.335 10.32 32.465 ;
		RECT	8.56 29.915 8.61 30.045 ;
		RECT	10.27 29.915 10.32 30.045 ;
		RECT	6.22 29.455 6.27 29.585 ;
		RECT	7.5 29.455 7.55 29.585 ;
		RECT	9.04 29.455 9.09 29.585 ;
		RECT	9.315 29.455 9.365 29.585 ;
		RECT	9.72 29.455 9.77 29.585 ;
		RECT	11.025 29.455 11.075 29.585 ;
		RECT	12.79 29.455 12.84 29.585 ;
		RECT	6.225 27.035 6.275 27.165 ;
		RECT	7.5 27.035 7.55 27.165 ;
		RECT	9.04 27.035 9.09 27.165 ;
		RECT	9.315 27.035 9.365 27.165 ;
		RECT	11.025 27.035 11.075 27.165 ;
		RECT	12.79 27.035 12.84 27.165 ;
		RECT	7.18 26.805 7.23 26.935 ;
		RECT	14.14 26.805 14.19 26.935 ;
		RECT	8.56 29.455 8.61 29.585 ;
		RECT	10.27 29.455 10.32 29.585 ;
		RECT	8.56 27.035 8.61 27.165 ;
		RECT	10.27 27.035 10.32 27.165 ;
		RECT	6.22 26.575 6.27 26.705 ;
		RECT	7.5 26.575 7.55 26.705 ;
		RECT	9.04 26.575 9.09 26.705 ;
		RECT	9.315 26.575 9.365 26.705 ;
		RECT	9.72 26.575 9.77 26.705 ;
		RECT	11.025 26.575 11.075 26.705 ;
		RECT	12.79 26.575 12.84 26.705 ;
		RECT	6.225 24.155 6.275 24.285 ;
		RECT	7.5 24.155 7.55 24.285 ;
		RECT	9.04 24.155 9.09 24.285 ;
		RECT	9.315 24.155 9.365 24.285 ;
		RECT	11.025 24.155 11.075 24.285 ;
		RECT	12.79 24.155 12.84 24.285 ;
		RECT	7.18 23.925 7.23 24.055 ;
		RECT	14.14 23.925 14.19 24.055 ;
		RECT	8.56 26.575 8.61 26.705 ;
		RECT	10.27 26.575 10.32 26.705 ;
		RECT	8.56 24.155 8.61 24.285 ;
		RECT	10.27 24.155 10.32 24.285 ;
		RECT	6.22 23.695 6.27 23.825 ;
		RECT	7.5 23.695 7.55 23.825 ;
		RECT	9.04 23.695 9.09 23.825 ;
		RECT	9.315 23.695 9.365 23.825 ;
		RECT	9.72 23.695 9.77 23.825 ;
		RECT	11.025 23.695 11.075 23.825 ;
		RECT	12.79 23.695 12.84 23.825 ;
		RECT	6.225 21.275 6.275 21.405 ;
		RECT	7.5 21.275 7.55 21.405 ;
		RECT	9.04 21.275 9.09 21.405 ;
		RECT	9.315 21.275 9.365 21.405 ;
		RECT	11.025 21.275 11.075 21.405 ;
		RECT	12.79 21.275 12.84 21.405 ;
		RECT	7.18 21.045 7.23 21.175 ;
		RECT	14.14 21.045 14.19 21.175 ;
		RECT	8.56 23.695 8.61 23.825 ;
		RECT	10.27 23.695 10.32 23.825 ;
		RECT	8.56 21.275 8.61 21.405 ;
		RECT	10.27 21.275 10.32 21.405 ;
		RECT	6.22 20.815 6.27 20.945 ;
		RECT	7.5 20.815 7.55 20.945 ;
		RECT	9.04 20.815 9.09 20.945 ;
		RECT	9.315 20.815 9.365 20.945 ;
		RECT	9.72 20.815 9.77 20.945 ;
		RECT	11.025 20.815 11.075 20.945 ;
		RECT	12.79 20.815 12.84 20.945 ;
		RECT	6.225 18.395 6.275 18.525 ;
		RECT	7.5 18.395 7.55 18.525 ;
		RECT	9.04 18.395 9.09 18.525 ;
		RECT	9.315 18.395 9.365 18.525 ;
		RECT	11.025 18.395 11.075 18.525 ;
		RECT	12.79 18.395 12.84 18.525 ;
		RECT	7.18 18.165 7.23 18.295 ;
		RECT	14.14 18.165 14.19 18.295 ;
		RECT	8.56 20.815 8.61 20.945 ;
		RECT	10.27 20.815 10.32 20.945 ;
		RECT	8.56 18.395 8.61 18.525 ;
		RECT	10.27 18.395 10.32 18.525 ;
		RECT	6.22 17.935 6.27 18.065 ;
		RECT	7.5 17.935 7.55 18.065 ;
		RECT	9.04 17.935 9.09 18.065 ;
		RECT	9.315 17.935 9.365 18.065 ;
		RECT	9.72 17.935 9.77 18.065 ;
		RECT	11.025 17.935 11.075 18.065 ;
		RECT	12.79 17.935 12.84 18.065 ;
		RECT	6.225 15.515 6.275 15.645 ;
		RECT	7.5 15.515 7.55 15.645 ;
		RECT	9.04 15.515 9.09 15.645 ;
		RECT	9.315 15.515 9.365 15.645 ;
		RECT	11.025 15.515 11.075 15.645 ;
		RECT	12.79 15.515 12.84 15.645 ;
		RECT	7.18 15.285 7.23 15.415 ;
		RECT	14.14 15.285 14.19 15.415 ;
		RECT	8.56 17.935 8.61 18.065 ;
		RECT	10.27 17.935 10.32 18.065 ;
		RECT	8.56 15.515 8.61 15.645 ;
		RECT	10.27 15.515 10.32 15.645 ;
		RECT	6.22 15.055 6.27 15.185 ;
		RECT	7.5 15.055 7.55 15.185 ;
		RECT	9.04 15.055 9.09 15.185 ;
		RECT	9.315 15.055 9.365 15.185 ;
		RECT	9.72 15.055 9.77 15.185 ;
		RECT	11.025 15.055 11.075 15.185 ;
		RECT	12.79 15.055 12.84 15.185 ;
		RECT	6.225 12.635 6.275 12.765 ;
		RECT	7.5 12.635 7.55 12.765 ;
		RECT	9.04 12.635 9.09 12.765 ;
		RECT	9.315 12.635 9.365 12.765 ;
		RECT	11.025 12.635 11.075 12.765 ;
		RECT	12.79 12.635 12.84 12.765 ;
		RECT	7.18 12.405 7.23 12.535 ;
		RECT	14.14 12.405 14.19 12.535 ;
		RECT	8.56 15.055 8.61 15.185 ;
		RECT	10.27 15.055 10.32 15.185 ;
		RECT	8.56 12.635 8.61 12.765 ;
		RECT	10.27 12.635 10.32 12.765 ;
		RECT	6.22 12.175 6.27 12.305 ;
		RECT	7.5 12.175 7.55 12.305 ;
		RECT	9.04 12.175 9.09 12.305 ;
		RECT	9.315 12.175 9.365 12.305 ;
		RECT	9.72 12.175 9.77 12.305 ;
		RECT	11.025 12.175 11.075 12.305 ;
		RECT	12.79 12.175 12.84 12.305 ;
		RECT	6.225 9.755 6.275 9.885 ;
		RECT	7.5 9.755 7.55 9.885 ;
		RECT	9.04 9.755 9.09 9.885 ;
		RECT	9.315 9.755 9.365 9.885 ;
		RECT	11.025 9.755 11.075 9.885 ;
		RECT	12.79 9.755 12.84 9.885 ;
		RECT	7.18 9.525 7.23 9.655 ;
		RECT	14.14 9.525 14.19 9.655 ;
		RECT	8.56 12.175 8.61 12.305 ;
		RECT	10.27 12.175 10.32 12.305 ;
		RECT	8.56 9.755 8.61 9.885 ;
		RECT	10.27 9.755 10.32 9.885 ;
		RECT	6.22 9.295 6.27 9.425 ;
		RECT	7.5 9.295 7.55 9.425 ;
		RECT	9.04 9.295 9.09 9.425 ;
		RECT	9.315 9.295 9.365 9.425 ;
		RECT	9.72 9.295 9.77 9.425 ;
		RECT	11.025 9.295 11.075 9.425 ;
		RECT	12.79 9.295 12.84 9.425 ;
		RECT	6.225 6.875 6.275 7.005 ;
		RECT	7.5 6.875 7.55 7.005 ;
		RECT	9.04 6.875 9.09 7.005 ;
		RECT	9.315 6.875 9.365 7.005 ;
		RECT	11.025 6.875 11.075 7.005 ;
		RECT	12.79 6.875 12.84 7.005 ;
		RECT	7.18 6.645 7.23 6.775 ;
		RECT	14.14 6.645 14.19 6.775 ;
		RECT	8.56 9.295 8.61 9.425 ;
		RECT	10.27 9.295 10.32 9.425 ;
		RECT	8.56 6.875 8.61 7.005 ;
		RECT	10.27 6.875 10.32 7.005 ;
		RECT	6.22 6.415 6.27 6.545 ;
		RECT	7.5 6.415 7.55 6.545 ;
		RECT	9.04 6.415 9.09 6.545 ;
		RECT	9.315 6.415 9.365 6.545 ;
		RECT	9.72 6.415 9.77 6.545 ;
		RECT	11.025 6.415 11.075 6.545 ;
		RECT	12.79 6.415 12.84 6.545 ;
		RECT	6.225 3.995 6.275 4.125 ;
		RECT	7.5 3.995 7.55 4.125 ;
		RECT	9.04 3.995 9.09 4.125 ;
		RECT	9.315 3.995 9.365 4.125 ;
		RECT	11.025 3.995 11.075 4.125 ;
		RECT	12.79 3.995 12.84 4.125 ;
		RECT	7.18 3.765 7.23 3.895 ;
		RECT	14.14 3.765 14.19 3.895 ;
		RECT	8.56 6.415 8.61 6.545 ;
		RECT	10.27 6.415 10.32 6.545 ;
		RECT	8.56 3.995 8.61 4.125 ;
		RECT	10.27 3.995 10.32 4.125 ;
		RECT	6.22 3.535 6.27 3.665 ;
		RECT	7.5 3.535 7.55 3.665 ;
		RECT	9.04 3.535 9.09 3.665 ;
		RECT	9.315 3.535 9.365 3.665 ;
		RECT	9.72 3.535 9.77 3.665 ;
		RECT	11.025 3.535 11.075 3.665 ;
		RECT	12.79 3.535 12.84 3.665 ;
		RECT	6.225 1.115 6.275 1.245 ;
		RECT	7.5 1.115 7.55 1.245 ;
		RECT	9.04 1.115 9.09 1.245 ;
		RECT	9.315 1.115 9.365 1.245 ;
		RECT	11.025 1.115 11.075 1.245 ;
		RECT	12.79 1.115 12.84 1.245 ;
		RECT	7.18 0.885 7.23 1.015 ;
		RECT	14.14 0.885 14.19 1.015 ;
		RECT	8.56 3.535 8.61 3.665 ;
		RECT	10.27 3.535 10.32 3.665 ;
		RECT	8.56 1.115 8.61 1.245 ;
		RECT	10.27 1.115 10.32 1.245 ;
		RECT	6.22 184.975 6.27 185.105 ;
		RECT	7.5 184.975 7.55 185.105 ;
		RECT	9.04 184.975 9.09 185.105 ;
		RECT	9.315 184.975 9.365 185.105 ;
		RECT	9.72 184.975 9.77 185.105 ;
		RECT	11.025 184.975 11.075 185.105 ;
		RECT	12.79 184.975 12.84 185.105 ;
		RECT	6.225 182.555 6.275 182.685 ;
		RECT	7.5 182.555 7.55 182.685 ;
		RECT	9.04 182.555 9.09 182.685 ;
		RECT	9.315 182.555 9.365 182.685 ;
		RECT	11.025 182.555 11.075 182.685 ;
		RECT	12.79 182.555 12.84 182.685 ;
		RECT	7.18 182.325 7.23 182.455 ;
		RECT	14.14 182.325 14.19 182.455 ;
		RECT	8.56 184.975 8.61 185.105 ;
		RECT	10.27 184.975 10.32 185.105 ;
		RECT	8.56 182.555 8.61 182.685 ;
		RECT	10.27 182.555 10.32 182.685 ;
		RECT	6.22 182.095 6.27 182.225 ;
		RECT	7.5 182.095 7.55 182.225 ;
		RECT	9.04 182.095 9.09 182.225 ;
		RECT	9.315 182.095 9.365 182.225 ;
		RECT	9.72 182.095 9.77 182.225 ;
		RECT	11.025 182.095 11.075 182.225 ;
		RECT	12.79 182.095 12.84 182.225 ;
		RECT	6.225 179.675 6.275 179.805 ;
		RECT	7.5 179.675 7.55 179.805 ;
		RECT	9.04 179.675 9.09 179.805 ;
		RECT	9.315 179.675 9.365 179.805 ;
		RECT	11.025 179.675 11.075 179.805 ;
		RECT	12.79 179.675 12.84 179.805 ;
		RECT	7.18 179.445 7.23 179.575 ;
		RECT	14.14 179.445 14.19 179.575 ;
		RECT	8.56 182.095 8.61 182.225 ;
		RECT	10.27 182.095 10.32 182.225 ;
		RECT	8.56 179.675 8.61 179.805 ;
		RECT	10.27 179.675 10.32 179.805 ;
		RECT	6.22 179.215 6.27 179.345 ;
		RECT	7.5 179.215 7.55 179.345 ;
		RECT	9.04 179.215 9.09 179.345 ;
		RECT	9.315 179.215 9.365 179.345 ;
		RECT	9.72 179.215 9.77 179.345 ;
		RECT	11.025 179.215 11.075 179.345 ;
		RECT	12.79 179.215 12.84 179.345 ;
		RECT	6.225 176.795 6.275 176.925 ;
		RECT	7.5 176.795 7.55 176.925 ;
		RECT	9.04 176.795 9.09 176.925 ;
		RECT	9.315 176.795 9.365 176.925 ;
		RECT	11.025 176.795 11.075 176.925 ;
		RECT	12.79 176.795 12.84 176.925 ;
		RECT	7.18 176.565 7.23 176.695 ;
		RECT	14.14 176.565 14.19 176.695 ;
		RECT	8.56 179.215 8.61 179.345 ;
		RECT	10.27 179.215 10.32 179.345 ;
		RECT	8.56 176.795 8.61 176.925 ;
		RECT	10.27 176.795 10.32 176.925 ;
		RECT	6.22 176.335 6.27 176.465 ;
		RECT	7.5 176.335 7.55 176.465 ;
		RECT	9.04 176.335 9.09 176.465 ;
		RECT	9.315 176.335 9.365 176.465 ;
		RECT	9.72 176.335 9.77 176.465 ;
		RECT	11.025 176.335 11.075 176.465 ;
		RECT	12.79 176.335 12.84 176.465 ;
		RECT	6.225 173.915 6.275 174.045 ;
		RECT	7.5 173.915 7.55 174.045 ;
		RECT	9.04 173.915 9.09 174.045 ;
		RECT	9.315 173.915 9.365 174.045 ;
		RECT	11.025 173.915 11.075 174.045 ;
		RECT	12.79 173.915 12.84 174.045 ;
		RECT	7.18 173.685 7.23 173.815 ;
		RECT	14.14 173.685 14.19 173.815 ;
		RECT	8.56 176.335 8.61 176.465 ;
		RECT	10.27 176.335 10.32 176.465 ;
		RECT	8.56 173.915 8.61 174.045 ;
		RECT	10.27 173.915 10.32 174.045 ;
		RECT	6.22 173.455 6.27 173.585 ;
		RECT	7.5 173.455 7.55 173.585 ;
		RECT	9.04 173.455 9.09 173.585 ;
		RECT	9.315 173.455 9.365 173.585 ;
		RECT	9.72 173.455 9.77 173.585 ;
		RECT	11.025 173.455 11.075 173.585 ;
		RECT	12.79 173.455 12.84 173.585 ;
		RECT	6.225 171.035 6.275 171.165 ;
		RECT	7.5 171.035 7.55 171.165 ;
		RECT	9.04 171.035 9.09 171.165 ;
		RECT	9.315 171.035 9.365 171.165 ;
		RECT	11.025 171.035 11.075 171.165 ;
		RECT	12.79 171.035 12.84 171.165 ;
		RECT	7.18 170.805 7.23 170.935 ;
		RECT	14.14 170.805 14.19 170.935 ;
		RECT	8.56 173.455 8.61 173.585 ;
		RECT	10.27 173.455 10.32 173.585 ;
		RECT	8.56 171.035 8.61 171.165 ;
		RECT	10.27 171.035 10.32 171.165 ;
		RECT	6.22 170.575 6.27 170.705 ;
		RECT	7.5 170.575 7.55 170.705 ;
		RECT	9.04 170.575 9.09 170.705 ;
		RECT	9.315 170.575 9.365 170.705 ;
		RECT	9.72 170.575 9.77 170.705 ;
		RECT	11.025 170.575 11.075 170.705 ;
		RECT	12.79 170.575 12.84 170.705 ;
		RECT	6.225 168.155 6.275 168.285 ;
		RECT	7.5 168.155 7.55 168.285 ;
		RECT	9.04 168.155 9.09 168.285 ;
		RECT	9.315 168.155 9.365 168.285 ;
		RECT	11.025 168.155 11.075 168.285 ;
		RECT	12.79 168.155 12.84 168.285 ;
		RECT	7.18 167.925 7.23 168.055 ;
		RECT	14.14 167.925 14.19 168.055 ;
		RECT	8.56 170.575 8.61 170.705 ;
		RECT	10.27 170.575 10.32 170.705 ;
		RECT	8.56 168.155 8.61 168.285 ;
		RECT	10.27 168.155 10.32 168.285 ;
		RECT	6.22 167.695 6.27 167.825 ;
		RECT	7.5 167.695 7.55 167.825 ;
		RECT	9.04 167.695 9.09 167.825 ;
		RECT	9.315 167.695 9.365 167.825 ;
		RECT	9.72 167.695 9.77 167.825 ;
		RECT	11.025 167.695 11.075 167.825 ;
		RECT	12.79 167.695 12.84 167.825 ;
		RECT	6.225 165.275 6.275 165.405 ;
		RECT	7.5 165.275 7.55 165.405 ;
		RECT	9.04 165.275 9.09 165.405 ;
		RECT	9.315 165.275 9.365 165.405 ;
		RECT	11.025 165.275 11.075 165.405 ;
		RECT	12.79 165.275 12.84 165.405 ;
		RECT	7.18 165.045 7.23 165.175 ;
		RECT	14.14 165.045 14.19 165.175 ;
		RECT	8.56 167.695 8.61 167.825 ;
		RECT	10.27 167.695 10.32 167.825 ;
		RECT	8.56 165.275 8.61 165.405 ;
		RECT	10.27 165.275 10.32 165.405 ;
		RECT	6.22 164.815 6.27 164.945 ;
		RECT	7.5 164.815 7.55 164.945 ;
		RECT	9.04 164.815 9.09 164.945 ;
		RECT	9.315 164.815 9.365 164.945 ;
		RECT	9.72 164.815 9.77 164.945 ;
		RECT	11.025 164.815 11.075 164.945 ;
		RECT	12.79 164.815 12.84 164.945 ;
		RECT	6.225 162.395 6.275 162.525 ;
		RECT	7.5 162.395 7.55 162.525 ;
		RECT	9.04 162.395 9.09 162.525 ;
		RECT	9.315 162.395 9.365 162.525 ;
		RECT	11.025 162.395 11.075 162.525 ;
		RECT	12.79 162.395 12.84 162.525 ;
		RECT	7.18 162.165 7.23 162.295 ;
		RECT	14.14 162.165 14.19 162.295 ;
		RECT	8.56 164.815 8.61 164.945 ;
		RECT	10.27 164.815 10.32 164.945 ;
		RECT	8.56 162.395 8.61 162.525 ;
		RECT	10.27 162.395 10.32 162.525 ;
		RECT	6.22 161.935 6.27 162.065 ;
		RECT	7.5 161.935 7.55 162.065 ;
		RECT	9.04 161.935 9.09 162.065 ;
		RECT	9.315 161.935 9.365 162.065 ;
		RECT	9.72 161.935 9.77 162.065 ;
		RECT	11.025 161.935 11.075 162.065 ;
		RECT	12.79 161.935 12.84 162.065 ;
		RECT	6.225 159.515 6.275 159.645 ;
		RECT	7.5 159.515 7.55 159.645 ;
		RECT	9.04 159.515 9.09 159.645 ;
		RECT	9.315 159.515 9.365 159.645 ;
		RECT	11.025 159.515 11.075 159.645 ;
		RECT	12.79 159.515 12.84 159.645 ;
		RECT	7.18 159.285 7.23 159.415 ;
		RECT	14.14 159.285 14.19 159.415 ;
		RECT	8.56 161.935 8.61 162.065 ;
		RECT	10.27 161.935 10.32 162.065 ;
		RECT	8.56 159.515 8.61 159.645 ;
		RECT	10.27 159.515 10.32 159.645 ;
		RECT	6.22 159.055 6.27 159.185 ;
		RECT	7.5 159.055 7.55 159.185 ;
		RECT	9.04 159.055 9.09 159.185 ;
		RECT	9.315 159.055 9.365 159.185 ;
		RECT	9.72 159.055 9.77 159.185 ;
		RECT	11.025 159.055 11.075 159.185 ;
		RECT	12.79 159.055 12.84 159.185 ;
		RECT	6.225 156.635 6.275 156.765 ;
		RECT	7.5 156.635 7.55 156.765 ;
		RECT	9.04 156.635 9.09 156.765 ;
		RECT	9.315 156.635 9.365 156.765 ;
		RECT	11.025 156.635 11.075 156.765 ;
		RECT	12.79 156.635 12.84 156.765 ;
		RECT	7.18 156.405 7.23 156.535 ;
		RECT	14.14 156.405 14.19 156.535 ;
		RECT	8.56 159.055 8.61 159.185 ;
		RECT	10.27 159.055 10.32 159.185 ;
		RECT	8.56 156.635 8.61 156.765 ;
		RECT	10.27 156.635 10.32 156.765 ;
		RECT	6.22 156.175 6.27 156.305 ;
		RECT	7.5 156.175 7.55 156.305 ;
		RECT	9.04 156.175 9.09 156.305 ;
		RECT	9.315 156.175 9.365 156.305 ;
		RECT	9.72 156.175 9.77 156.305 ;
		RECT	11.025 156.175 11.075 156.305 ;
		RECT	12.79 156.175 12.84 156.305 ;
		RECT	6.225 153.755 6.275 153.885 ;
		RECT	7.5 153.755 7.55 153.885 ;
		RECT	9.04 153.755 9.09 153.885 ;
		RECT	9.315 153.755 9.365 153.885 ;
		RECT	11.025 153.755 11.075 153.885 ;
		RECT	12.79 153.755 12.84 153.885 ;
		RECT	7.18 153.525 7.23 153.655 ;
		RECT	14.14 153.525 14.19 153.655 ;
		RECT	8.56 156.175 8.61 156.305 ;
		RECT	10.27 156.175 10.32 156.305 ;
		RECT	8.56 153.755 8.61 153.885 ;
		RECT	10.27 153.755 10.32 153.885 ;
		RECT	6.22 153.295 6.27 153.425 ;
		RECT	7.5 153.295 7.55 153.425 ;
		RECT	9.04 153.295 9.09 153.425 ;
		RECT	9.315 153.295 9.365 153.425 ;
		RECT	9.72 153.295 9.77 153.425 ;
		RECT	11.025 153.295 11.075 153.425 ;
		RECT	12.79 153.295 12.84 153.425 ;
		RECT	6.225 150.875 6.275 151.005 ;
		RECT	7.5 150.875 7.55 151.005 ;
		RECT	9.04 150.875 9.09 151.005 ;
		RECT	9.315 150.875 9.365 151.005 ;
		RECT	11.025 150.875 11.075 151.005 ;
		RECT	12.79 150.875 12.84 151.005 ;
		RECT	7.18 150.645 7.23 150.775 ;
		RECT	14.14 150.645 14.19 150.775 ;
		RECT	8.56 153.295 8.61 153.425 ;
		RECT	10.27 153.295 10.32 153.425 ;
		RECT	8.56 150.875 8.61 151.005 ;
		RECT	10.27 150.875 10.32 151.005 ;
		RECT	6.22 150.415 6.27 150.545 ;
		RECT	7.5 150.415 7.55 150.545 ;
		RECT	9.04 150.415 9.09 150.545 ;
		RECT	9.315 150.415 9.365 150.545 ;
		RECT	9.72 150.415 9.77 150.545 ;
		RECT	11.025 150.415 11.075 150.545 ;
		RECT	12.79 150.415 12.84 150.545 ;
		RECT	6.225 147.995 6.275 148.125 ;
		RECT	7.5 147.995 7.55 148.125 ;
		RECT	9.04 147.995 9.09 148.125 ;
		RECT	9.315 147.995 9.365 148.125 ;
		RECT	11.025 147.995 11.075 148.125 ;
		RECT	12.79 147.995 12.84 148.125 ;
		RECT	7.18 147.765 7.23 147.895 ;
		RECT	14.14 147.765 14.19 147.895 ;
		RECT	8.56 150.415 8.61 150.545 ;
		RECT	10.27 150.415 10.32 150.545 ;
		RECT	8.56 147.995 8.61 148.125 ;
		RECT	10.27 147.995 10.32 148.125 ;
		RECT	6.22 147.535 6.27 147.665 ;
		RECT	7.5 147.535 7.55 147.665 ;
		RECT	9.04 147.535 9.09 147.665 ;
		RECT	9.315 147.535 9.365 147.665 ;
		RECT	9.72 147.535 9.77 147.665 ;
		RECT	11.025 147.535 11.075 147.665 ;
		RECT	12.79 147.535 12.84 147.665 ;
		RECT	6.225 145.115 6.275 145.245 ;
		RECT	7.5 145.115 7.55 145.245 ;
		RECT	9.04 145.115 9.09 145.245 ;
		RECT	9.315 145.115 9.365 145.245 ;
		RECT	11.025 145.115 11.075 145.245 ;
		RECT	12.79 145.115 12.84 145.245 ;
		RECT	7.18 144.885 7.23 145.015 ;
		RECT	14.14 144.885 14.19 145.015 ;
		RECT	8.56 147.535 8.61 147.665 ;
		RECT	10.27 147.535 10.32 147.665 ;
		RECT	8.56 145.115 8.61 145.245 ;
		RECT	10.27 145.115 10.32 145.245 ;
		RECT	6.22 144.655 6.27 144.785 ;
		RECT	7.5 144.655 7.55 144.785 ;
		RECT	9.04 144.655 9.09 144.785 ;
		RECT	9.315 144.655 9.365 144.785 ;
		RECT	9.72 144.655 9.77 144.785 ;
		RECT	11.025 144.655 11.075 144.785 ;
		RECT	12.79 144.655 12.84 144.785 ;
		RECT	6.225 142.235 6.275 142.365 ;
		RECT	7.5 142.235 7.55 142.365 ;
		RECT	9.04 142.235 9.09 142.365 ;
		RECT	9.315 142.235 9.365 142.365 ;
		RECT	11.025 142.235 11.075 142.365 ;
		RECT	12.79 142.235 12.84 142.365 ;
		RECT	7.18 142.005 7.23 142.135 ;
		RECT	14.14 142.005 14.19 142.135 ;
		RECT	8.56 144.655 8.61 144.785 ;
		RECT	10.27 144.655 10.32 144.785 ;
		RECT	8.56 142.235 8.61 142.365 ;
		RECT	10.27 142.235 10.32 142.365 ;
		RECT	6.22 141.775 6.27 141.905 ;
		RECT	7.5 141.775 7.55 141.905 ;
		RECT	9.04 141.775 9.09 141.905 ;
		RECT	9.315 141.775 9.365 141.905 ;
		RECT	9.72 141.775 9.77 141.905 ;
		RECT	11.025 141.775 11.075 141.905 ;
		RECT	12.79 141.775 12.84 141.905 ;
		RECT	6.225 139.355 6.275 139.485 ;
		RECT	7.5 139.355 7.55 139.485 ;
		RECT	9.04 139.355 9.09 139.485 ;
		RECT	9.315 139.355 9.365 139.485 ;
		RECT	11.025 139.355 11.075 139.485 ;
		RECT	12.79 139.355 12.84 139.485 ;
		RECT	7.18 139.125 7.23 139.255 ;
		RECT	14.14 139.125 14.19 139.255 ;
		RECT	8.56 141.775 8.61 141.905 ;
		RECT	10.27 141.775 10.32 141.905 ;
		RECT	8.56 139.355 8.61 139.485 ;
		RECT	10.27 139.355 10.32 139.485 ;
		RECT	6.22 138.895 6.27 139.025 ;
		RECT	7.5 138.895 7.55 139.025 ;
		RECT	9.04 138.895 9.09 139.025 ;
		RECT	9.315 138.895 9.365 139.025 ;
		RECT	9.72 138.895 9.77 139.025 ;
		RECT	11.025 138.895 11.075 139.025 ;
		RECT	12.79 138.895 12.84 139.025 ;
		RECT	6.225 136.475 6.275 136.605 ;
		RECT	7.5 136.475 7.55 136.605 ;
		RECT	9.04 136.475 9.09 136.605 ;
		RECT	9.315 136.475 9.365 136.605 ;
		RECT	11.025 136.475 11.075 136.605 ;
		RECT	12.79 136.475 12.84 136.605 ;
		RECT	7.18 136.245 7.23 136.375 ;
		RECT	14.14 136.245 14.19 136.375 ;
		RECT	8.56 138.895 8.61 139.025 ;
		RECT	10.27 138.895 10.32 139.025 ;
		RECT	8.56 136.475 8.61 136.605 ;
		RECT	10.27 136.475 10.32 136.605 ;
		RECT	6.22 136.015 6.27 136.145 ;
		RECT	7.5 136.015 7.55 136.145 ;
		RECT	9.04 136.015 9.09 136.145 ;
		RECT	9.315 136.015 9.365 136.145 ;
		RECT	9.72 136.015 9.77 136.145 ;
		RECT	11.025 136.015 11.075 136.145 ;
		RECT	12.79 136.015 12.84 136.145 ;
		RECT	6.225 133.595 6.275 133.725 ;
		RECT	7.5 133.595 7.55 133.725 ;
		RECT	9.04 133.595 9.09 133.725 ;
		RECT	9.315 133.595 9.365 133.725 ;
		RECT	11.025 133.595 11.075 133.725 ;
		RECT	12.79 133.595 12.84 133.725 ;
		RECT	7.18 133.365 7.23 133.495 ;
		RECT	14.14 133.365 14.19 133.495 ;
		RECT	8.56 136.015 8.61 136.145 ;
		RECT	10.27 136.015 10.32 136.145 ;
		RECT	8.56 133.595 8.61 133.725 ;
		RECT	10.27 133.595 10.32 133.725 ;
		RECT	6.22 133.135 6.27 133.265 ;
		RECT	7.5 133.135 7.55 133.265 ;
		RECT	9.04 133.135 9.09 133.265 ;
		RECT	9.315 133.135 9.365 133.265 ;
		RECT	9.72 133.135 9.77 133.265 ;
		RECT	11.025 133.135 11.075 133.265 ;
		RECT	12.79 133.135 12.84 133.265 ;
		RECT	6.225 130.715 6.275 130.845 ;
		RECT	7.5 130.715 7.55 130.845 ;
		RECT	9.04 130.715 9.09 130.845 ;
		RECT	9.315 130.715 9.365 130.845 ;
		RECT	11.025 130.715 11.075 130.845 ;
		RECT	12.79 130.715 12.84 130.845 ;
		RECT	7.18 130.485 7.23 130.615 ;
		RECT	14.14 130.485 14.19 130.615 ;
		RECT	8.56 133.135 8.61 133.265 ;
		RECT	10.27 133.135 10.32 133.265 ;
		RECT	8.56 130.715 8.61 130.845 ;
		RECT	10.27 130.715 10.32 130.845 ;
		RECT	6.22 130.255 6.27 130.385 ;
		RECT	7.5 130.255 7.55 130.385 ;
		RECT	9.04 130.255 9.09 130.385 ;
		RECT	9.315 130.255 9.365 130.385 ;
		RECT	9.72 130.255 9.77 130.385 ;
		RECT	11.025 130.255 11.075 130.385 ;
		RECT	12.79 130.255 12.84 130.385 ;
		RECT	6.225 127.835 6.275 127.965 ;
		RECT	7.5 127.835 7.55 127.965 ;
		RECT	9.04 127.835 9.09 127.965 ;
		RECT	9.315 127.835 9.365 127.965 ;
		RECT	11.025 127.835 11.075 127.965 ;
		RECT	12.79 127.835 12.84 127.965 ;
		RECT	7.18 127.605 7.23 127.735 ;
		RECT	14.14 127.605 14.19 127.735 ;
		RECT	8.56 130.255 8.61 130.385 ;
		RECT	10.27 130.255 10.32 130.385 ;
		RECT	8.56 127.835 8.61 127.965 ;
		RECT	10.27 127.835 10.32 127.965 ;
		RECT	6.22 127.375 6.27 127.505 ;
		RECT	7.5 127.375 7.55 127.505 ;
		RECT	9.04 127.375 9.09 127.505 ;
		RECT	9.315 127.375 9.365 127.505 ;
		RECT	9.72 127.375 9.77 127.505 ;
		RECT	11.025 127.375 11.075 127.505 ;
		RECT	12.79 127.375 12.84 127.505 ;
		RECT	14.33 182.095 14.38 182.225 ;
		RECT	6.22 181.635 6.27 181.765 ;
		RECT	7.5 181.635 7.55 181.765 ;
		RECT	9.04 181.635 9.09 181.765 ;
		RECT	9.315 181.635 9.365 181.765 ;
		RECT	9.72 181.635 9.77 181.765 ;
		RECT	11.025 181.635 11.075 181.765 ;
		RECT	12.79 181.635 12.84 181.765 ;
		RECT	14.33 179.675 14.38 179.805 ;
		RECT	5.675 179.445 5.725 179.575 ;
		RECT	6.065 179.445 6.115 179.575 ;
		RECT	6.725 179.445 6.775 179.575 ;
		RECT	8.42 179.445 8.47 179.575 ;
		RECT	8.77 179.445 8.82 179.575 ;
		RECT	11.555 179.445 11.605 179.575 ;
		RECT	11.815 179.445 11.865 179.575 ;
		RECT	12.52 179.445 12.57 179.575 ;
		RECT	13.98 179.445 14.03 179.575 ;
		RECT	14.33 156.175 14.38 156.305 ;
		RECT	6.22 155.715 6.27 155.845 ;
		RECT	7.5 155.715 7.55 155.845 ;
		RECT	9.04 155.715 9.09 155.845 ;
		RECT	9.315 155.715 9.365 155.845 ;
		RECT	9.72 155.715 9.77 155.845 ;
		RECT	11.025 155.715 11.075 155.845 ;
		RECT	12.79 155.715 12.84 155.845 ;
		RECT	14.33 153.755 14.38 153.885 ;
		RECT	5.675 153.525 5.725 153.655 ;
		RECT	6.065 153.525 6.115 153.655 ;
		RECT	6.725 153.525 6.775 153.655 ;
		RECT	8.42 153.525 8.47 153.655 ;
		RECT	8.77 153.525 8.82 153.655 ;
		RECT	11.555 153.525 11.605 153.655 ;
		RECT	11.815 153.525 11.865 153.655 ;
		RECT	12.52 153.525 12.57 153.655 ;
		RECT	13.98 153.525 14.03 153.655 ;
		RECT	14.33 153.295 14.38 153.425 ;
		RECT	6.22 152.835 6.27 152.965 ;
		RECT	7.5 152.835 7.55 152.965 ;
		RECT	9.04 152.835 9.09 152.965 ;
		RECT	9.315 152.835 9.365 152.965 ;
		RECT	9.72 152.835 9.77 152.965 ;
		RECT	11.025 152.835 11.075 152.965 ;
		RECT	12.79 152.835 12.84 152.965 ;
		RECT	14.33 150.875 14.38 151.005 ;
		RECT	5.675 150.645 5.725 150.775 ;
		RECT	6.065 150.645 6.115 150.775 ;
		RECT	6.725 150.645 6.775 150.775 ;
		RECT	8.42 150.645 8.47 150.775 ;
		RECT	8.77 150.645 8.82 150.775 ;
		RECT	11.555 150.645 11.605 150.775 ;
		RECT	11.815 150.645 11.865 150.775 ;
		RECT	12.52 150.645 12.57 150.775 ;
		RECT	13.98 150.645 14.03 150.775 ;
		RECT	14.33 150.415 14.38 150.545 ;
		RECT	6.22 149.955 6.27 150.085 ;
		RECT	7.5 149.955 7.55 150.085 ;
		RECT	9.04 149.955 9.09 150.085 ;
		RECT	9.315 149.955 9.365 150.085 ;
		RECT	9.72 149.955 9.77 150.085 ;
		RECT	11.025 149.955 11.075 150.085 ;
		RECT	12.79 149.955 12.84 150.085 ;
		RECT	14.33 147.995 14.38 148.125 ;
		RECT	5.675 147.765 5.725 147.895 ;
		RECT	6.065 147.765 6.115 147.895 ;
		RECT	6.725 147.765 6.775 147.895 ;
		RECT	8.42 147.765 8.47 147.895 ;
		RECT	8.77 147.765 8.82 147.895 ;
		RECT	11.555 147.765 11.605 147.895 ;
		RECT	11.815 147.765 11.865 147.895 ;
		RECT	12.52 147.765 12.57 147.895 ;
		RECT	13.98 147.765 14.03 147.895 ;
		RECT	14.33 147.535 14.38 147.665 ;
		RECT	6.22 147.075 6.27 147.205 ;
		RECT	7.5 147.075 7.55 147.205 ;
		RECT	9.04 147.075 9.09 147.205 ;
		RECT	9.315 147.075 9.365 147.205 ;
		RECT	9.72 147.075 9.77 147.205 ;
		RECT	11.025 147.075 11.075 147.205 ;
		RECT	12.79 147.075 12.84 147.205 ;
		RECT	14.33 145.115 14.38 145.245 ;
		RECT	5.675 144.885 5.725 145.015 ;
		RECT	6.065 144.885 6.115 145.015 ;
		RECT	6.725 144.885 6.775 145.015 ;
		RECT	8.42 144.885 8.47 145.015 ;
		RECT	8.77 144.885 8.82 145.015 ;
		RECT	11.555 144.885 11.605 145.015 ;
		RECT	11.815 144.885 11.865 145.015 ;
		RECT	12.52 144.885 12.57 145.015 ;
		RECT	13.98 144.885 14.03 145.015 ;
		RECT	14.33 144.655 14.38 144.785 ;
		RECT	6.22 144.195 6.27 144.325 ;
		RECT	7.5 144.195 7.55 144.325 ;
		RECT	9.04 144.195 9.09 144.325 ;
		RECT	9.315 144.195 9.365 144.325 ;
		RECT	9.72 144.195 9.77 144.325 ;
		RECT	11.025 144.195 11.075 144.325 ;
		RECT	12.79 144.195 12.84 144.325 ;
		RECT	14.33 142.235 14.38 142.365 ;
		RECT	5.675 142.005 5.725 142.135 ;
		RECT	6.065 142.005 6.115 142.135 ;
		RECT	6.725 142.005 6.775 142.135 ;
		RECT	8.42 142.005 8.47 142.135 ;
		RECT	8.77 142.005 8.82 142.135 ;
		RECT	11.555 142.005 11.605 142.135 ;
		RECT	11.815 142.005 11.865 142.135 ;
		RECT	12.52 142.005 12.57 142.135 ;
		RECT	13.98 142.005 14.03 142.135 ;
		RECT	14.33 141.775 14.38 141.905 ;
		RECT	6.22 141.315 6.27 141.445 ;
		RECT	7.5 141.315 7.55 141.445 ;
		RECT	9.04 141.315 9.09 141.445 ;
		RECT	9.315 141.315 9.365 141.445 ;
		RECT	9.72 141.315 9.77 141.445 ;
		RECT	11.025 141.315 11.075 141.445 ;
		RECT	12.79 141.315 12.84 141.445 ;
		RECT	14.33 139.355 14.38 139.485 ;
		RECT	5.675 139.125 5.725 139.255 ;
		RECT	6.065 139.125 6.115 139.255 ;
		RECT	6.725 139.125 6.775 139.255 ;
		RECT	8.42 139.125 8.47 139.255 ;
		RECT	8.77 139.125 8.82 139.255 ;
		RECT	11.555 139.125 11.605 139.255 ;
		RECT	11.815 139.125 11.865 139.255 ;
		RECT	12.52 139.125 12.57 139.255 ;
		RECT	13.98 139.125 14.03 139.255 ;
		RECT	14.33 138.895 14.38 139.025 ;
		RECT	6.22 138.435 6.27 138.565 ;
		RECT	7.5 138.435 7.55 138.565 ;
		RECT	9.04 138.435 9.09 138.565 ;
		RECT	9.315 138.435 9.365 138.565 ;
		RECT	9.72 138.435 9.77 138.565 ;
		RECT	11.025 138.435 11.075 138.565 ;
		RECT	12.79 138.435 12.84 138.565 ;
		RECT	14.33 136.475 14.38 136.605 ;
		RECT	5.675 136.245 5.725 136.375 ;
		RECT	6.065 136.245 6.115 136.375 ;
		RECT	6.725 136.245 6.775 136.375 ;
		RECT	8.42 136.245 8.47 136.375 ;
		RECT	8.77 136.245 8.82 136.375 ;
		RECT	11.555 136.245 11.605 136.375 ;
		RECT	11.815 136.245 11.865 136.375 ;
		RECT	12.52 136.245 12.57 136.375 ;
		RECT	13.98 136.245 14.03 136.375 ;
		RECT	14.33 136.015 14.38 136.145 ;
		RECT	6.22 135.555 6.27 135.685 ;
		RECT	7.5 135.555 7.55 135.685 ;
		RECT	9.04 135.555 9.09 135.685 ;
		RECT	9.315 135.555 9.365 135.685 ;
		RECT	9.72 135.555 9.77 135.685 ;
		RECT	11.025 135.555 11.075 135.685 ;
		RECT	12.79 135.555 12.84 135.685 ;
		RECT	14.33 133.595 14.38 133.725 ;
		RECT	5.675 133.365 5.725 133.495 ;
		RECT	6.065 133.365 6.115 133.495 ;
		RECT	6.725 133.365 6.775 133.495 ;
		RECT	8.42 133.365 8.47 133.495 ;
		RECT	8.77 133.365 8.82 133.495 ;
		RECT	11.555 133.365 11.605 133.495 ;
		RECT	11.815 133.365 11.865 133.495 ;
		RECT	12.52 133.365 12.57 133.495 ;
		RECT	13.98 133.365 14.03 133.495 ;
		RECT	14.33 133.135 14.38 133.265 ;
		RECT	6.22 132.675 6.27 132.805 ;
		RECT	7.5 132.675 7.55 132.805 ;
		RECT	9.04 132.675 9.09 132.805 ;
		RECT	9.315 132.675 9.365 132.805 ;
		RECT	9.72 132.675 9.77 132.805 ;
		RECT	11.025 132.675 11.075 132.805 ;
		RECT	12.79 132.675 12.84 132.805 ;
		RECT	14.33 130.715 14.38 130.845 ;
		RECT	5.675 130.485 5.725 130.615 ;
		RECT	6.065 130.485 6.115 130.615 ;
		RECT	6.725 130.485 6.775 130.615 ;
		RECT	8.42 130.485 8.47 130.615 ;
		RECT	8.77 130.485 8.82 130.615 ;
		RECT	11.555 130.485 11.605 130.615 ;
		RECT	11.815 130.485 11.865 130.615 ;
		RECT	12.52 130.485 12.57 130.615 ;
		RECT	13.98 130.485 14.03 130.615 ;
		RECT	14.33 130.255 14.38 130.385 ;
		RECT	6.22 129.795 6.27 129.925 ;
		RECT	7.5 129.795 7.55 129.925 ;
		RECT	9.04 129.795 9.09 129.925 ;
		RECT	9.315 129.795 9.365 129.925 ;
		RECT	9.72 129.795 9.77 129.925 ;
		RECT	11.025 129.795 11.075 129.925 ;
		RECT	12.79 129.795 12.84 129.925 ;
		RECT	14.33 127.835 14.38 127.965 ;
		RECT	5.675 127.605 5.725 127.735 ;
		RECT	6.065 127.605 6.115 127.735 ;
		RECT	6.725 127.605 6.775 127.735 ;
		RECT	8.42 127.605 8.47 127.735 ;
		RECT	8.77 127.605 8.82 127.735 ;
		RECT	11.555 127.605 11.605 127.735 ;
		RECT	11.815 127.605 11.865 127.735 ;
		RECT	12.52 127.605 12.57 127.735 ;
		RECT	13.98 127.605 14.03 127.735 ;
		RECT	14.33 179.215 14.38 179.345 ;
		RECT	6.22 178.755 6.27 178.885 ;
		RECT	7.5 178.755 7.55 178.885 ;
		RECT	9.04 178.755 9.09 178.885 ;
		RECT	9.315 178.755 9.365 178.885 ;
		RECT	9.72 178.755 9.77 178.885 ;
		RECT	11.025 178.755 11.075 178.885 ;
		RECT	12.79 178.755 12.84 178.885 ;
		RECT	14.33 176.795 14.38 176.925 ;
		RECT	5.675 176.565 5.725 176.695 ;
		RECT	6.065 176.565 6.115 176.695 ;
		RECT	6.725 176.565 6.775 176.695 ;
		RECT	8.42 176.565 8.47 176.695 ;
		RECT	8.77 176.565 8.82 176.695 ;
		RECT	11.555 176.565 11.605 176.695 ;
		RECT	11.815 176.565 11.865 176.695 ;
		RECT	12.52 176.565 12.57 176.695 ;
		RECT	13.98 176.565 14.03 176.695 ;
		RECT	14.33 127.375 14.38 127.505 ;
		RECT	6.22 126.915 6.27 127.045 ;
		RECT	7.5 126.915 7.55 127.045 ;
		RECT	9.04 126.915 9.09 127.045 ;
		RECT	9.315 126.915 9.365 127.045 ;
		RECT	9.72 126.915 9.77 127.045 ;
		RECT	11.025 126.915 11.075 127.045 ;
		RECT	12.79 126.915 12.84 127.045 ;
		RECT	14.33 124.955 14.38 125.085 ;
		RECT	5.675 124.725 5.725 124.855 ;
		RECT	6.065 124.725 6.115 124.855 ;
		RECT	6.725 124.725 6.775 124.855 ;
		RECT	8.42 124.725 8.47 124.855 ;
		RECT	8.77 124.725 8.82 124.855 ;
		RECT	11.555 124.725 11.605 124.855 ;
		RECT	11.815 124.725 11.865 124.855 ;
		RECT	12.52 124.725 12.57 124.855 ;
		RECT	13.98 124.725 14.03 124.855 ;
		RECT	14.33 124.495 14.38 124.625 ;
		RECT	6.22 124.035 6.27 124.165 ;
		RECT	7.5 124.035 7.55 124.165 ;
		RECT	9.04 124.035 9.09 124.165 ;
		RECT	9.315 124.035 9.365 124.165 ;
		RECT	9.72 124.035 9.77 124.165 ;
		RECT	11.025 124.035 11.075 124.165 ;
		RECT	12.79 124.035 12.84 124.165 ;
		RECT	14.33 122.075 14.38 122.205 ;
		RECT	5.675 121.845 5.725 121.975 ;
		RECT	6.065 121.845 6.115 121.975 ;
		RECT	6.725 121.845 6.775 121.975 ;
		RECT	8.42 121.845 8.47 121.975 ;
		RECT	8.77 121.845 8.82 121.975 ;
		RECT	11.555 121.845 11.605 121.975 ;
		RECT	11.815 121.845 11.865 121.975 ;
		RECT	12.52 121.845 12.57 121.975 ;
		RECT	13.98 121.845 14.03 121.975 ;
		RECT	14.33 121.615 14.38 121.745 ;
		RECT	6.22 121.155 6.27 121.285 ;
		RECT	7.5 121.155 7.55 121.285 ;
		RECT	9.04 121.155 9.09 121.285 ;
		RECT	9.315 121.155 9.365 121.285 ;
		RECT	9.72 121.155 9.77 121.285 ;
		RECT	11.025 121.155 11.075 121.285 ;
		RECT	12.79 121.155 12.84 121.285 ;
		RECT	14.33 119.195 14.38 119.325 ;
		RECT	5.675 118.965 5.725 119.095 ;
		RECT	6.065 118.965 6.115 119.095 ;
		RECT	6.725 118.965 6.775 119.095 ;
		RECT	8.42 118.965 8.47 119.095 ;
		RECT	8.77 118.965 8.82 119.095 ;
		RECT	11.555 118.965 11.605 119.095 ;
		RECT	11.815 118.965 11.865 119.095 ;
		RECT	12.52 118.965 12.57 119.095 ;
		RECT	13.98 118.965 14.03 119.095 ;
		RECT	14.33 118.735 14.38 118.865 ;
		RECT	6.22 118.275 6.27 118.405 ;
		RECT	7.5 118.275 7.55 118.405 ;
		RECT	9.04 118.275 9.09 118.405 ;
		RECT	9.315 118.275 9.365 118.405 ;
		RECT	9.72 118.275 9.77 118.405 ;
		RECT	11.025 118.275 11.075 118.405 ;
		RECT	12.79 118.275 12.84 118.405 ;
		RECT	14.33 116.315 14.38 116.445 ;
		RECT	5.675 116.085 5.725 116.215 ;
		RECT	6.065 116.085 6.115 116.215 ;
		RECT	6.725 116.085 6.775 116.215 ;
		RECT	8.42 116.085 8.47 116.215 ;
		RECT	8.77 116.085 8.82 116.215 ;
		RECT	11.555 116.085 11.605 116.215 ;
		RECT	11.815 116.085 11.865 116.215 ;
		RECT	12.52 116.085 12.57 116.215 ;
		RECT	13.98 116.085 14.03 116.215 ;
		RECT	14.33 115.855 14.38 115.985 ;
		RECT	6.22 115.395 6.27 115.525 ;
		RECT	7.5 115.395 7.55 115.525 ;
		RECT	9.04 115.395 9.09 115.525 ;
		RECT	9.315 115.395 9.365 115.525 ;
		RECT	9.72 115.395 9.77 115.525 ;
		RECT	11.025 115.395 11.075 115.525 ;
		RECT	12.79 115.395 12.84 115.525 ;
		RECT	14.33 113.435 14.38 113.565 ;
		RECT	5.675 113.205 5.725 113.335 ;
		RECT	6.065 113.205 6.115 113.335 ;
		RECT	6.725 113.205 6.775 113.335 ;
		RECT	8.42 113.205 8.47 113.335 ;
		RECT	8.77 113.205 8.82 113.335 ;
		RECT	11.555 113.205 11.605 113.335 ;
		RECT	11.815 113.205 11.865 113.335 ;
		RECT	12.52 113.205 12.57 113.335 ;
		RECT	13.98 113.205 14.03 113.335 ;
		RECT	14.33 112.975 14.38 113.105 ;
		RECT	6.22 112.515 6.27 112.645 ;
		RECT	7.5 112.515 7.55 112.645 ;
		RECT	9.04 112.515 9.09 112.645 ;
		RECT	9.315 112.515 9.365 112.645 ;
		RECT	9.72 112.515 9.77 112.645 ;
		RECT	11.025 112.515 11.075 112.645 ;
		RECT	12.79 112.515 12.84 112.645 ;
		RECT	14.33 110.555 14.38 110.685 ;
		RECT	5.675 110.325 5.725 110.455 ;
		RECT	6.065 110.325 6.115 110.455 ;
		RECT	6.725 110.325 6.775 110.455 ;
		RECT	8.42 110.325 8.47 110.455 ;
		RECT	8.77 110.325 8.82 110.455 ;
		RECT	11.555 110.325 11.605 110.455 ;
		RECT	11.815 110.325 11.865 110.455 ;
		RECT	12.52 110.325 12.57 110.455 ;
		RECT	13.98 110.325 14.03 110.455 ;
		RECT	14.33 110.095 14.38 110.225 ;
		RECT	6.22 109.635 6.27 109.765 ;
		RECT	7.5 109.635 7.55 109.765 ;
		RECT	9.04 109.635 9.09 109.765 ;
		RECT	9.315 109.635 9.365 109.765 ;
		RECT	9.72 109.635 9.77 109.765 ;
		RECT	11.025 109.635 11.075 109.765 ;
		RECT	12.79 109.635 12.84 109.765 ;
		RECT	14.33 107.675 14.38 107.805 ;
		RECT	5.675 107.445 5.725 107.575 ;
		RECT	6.065 107.445 6.115 107.575 ;
		RECT	6.725 107.445 6.775 107.575 ;
		RECT	8.42 107.445 8.47 107.575 ;
		RECT	8.77 107.445 8.82 107.575 ;
		RECT	11.555 107.445 11.605 107.575 ;
		RECT	11.815 107.445 11.865 107.575 ;
		RECT	12.52 107.445 12.57 107.575 ;
		RECT	13.98 107.445 14.03 107.575 ;
		RECT	14.33 107.215 14.38 107.345 ;
		RECT	6.22 106.755 6.27 106.885 ;
		RECT	7.5 106.755 7.55 106.885 ;
		RECT	9.04 106.755 9.09 106.885 ;
		RECT	9.315 106.755 9.365 106.885 ;
		RECT	9.72 106.755 9.77 106.885 ;
		RECT	11.025 106.755 11.075 106.885 ;
		RECT	12.79 106.755 12.84 106.885 ;
		RECT	14.33 104.795 14.38 104.925 ;
		RECT	5.675 104.565 5.725 104.695 ;
		RECT	6.065 104.565 6.115 104.695 ;
		RECT	6.725 104.565 6.775 104.695 ;
		RECT	8.42 104.565 8.47 104.695 ;
		RECT	8.77 104.565 8.82 104.695 ;
		RECT	11.555 104.565 11.605 104.695 ;
		RECT	11.815 104.565 11.865 104.695 ;
		RECT	12.52 104.565 12.57 104.695 ;
		RECT	13.98 104.565 14.03 104.695 ;
		RECT	14.33 104.335 14.38 104.465 ;
		RECT	6.22 103.875 6.27 104.005 ;
		RECT	7.5 103.875 7.55 104.005 ;
		RECT	9.04 103.875 9.09 104.005 ;
		RECT	9.315 103.875 9.365 104.005 ;
		RECT	9.72 103.875 9.77 104.005 ;
		RECT	11.025 103.875 11.075 104.005 ;
		RECT	12.79 103.875 12.84 104.005 ;
		RECT	14.33 101.915 14.38 102.045 ;
		RECT	5.675 101.685 5.725 101.815 ;
		RECT	6.065 101.685 6.115 101.815 ;
		RECT	6.725 101.685 6.775 101.815 ;
		RECT	8.42 101.685 8.47 101.815 ;
		RECT	8.77 101.685 8.82 101.815 ;
		RECT	11.555 101.685 11.605 101.815 ;
		RECT	11.815 101.685 11.865 101.815 ;
		RECT	12.52 101.685 12.57 101.815 ;
		RECT	13.98 101.685 14.03 101.815 ;
		RECT	14.33 101.455 14.38 101.585 ;
		RECT	6.22 100.995 6.27 101.125 ;
		RECT	7.5 100.995 7.55 101.125 ;
		RECT	9.04 100.995 9.09 101.125 ;
		RECT	9.315 100.995 9.365 101.125 ;
		RECT	9.72 100.995 9.77 101.125 ;
		RECT	11.025 100.995 11.075 101.125 ;
		RECT	12.79 100.995 12.84 101.125 ;
		RECT	14.33 99.035 14.38 99.165 ;
		RECT	5.675 98.805 5.725 98.935 ;
		RECT	6.065 98.805 6.115 98.935 ;
		RECT	6.725 98.805 6.775 98.935 ;
		RECT	8.42 98.805 8.47 98.935 ;
		RECT	8.77 98.805 8.82 98.935 ;
		RECT	11.555 98.805 11.605 98.935 ;
		RECT	11.815 98.805 11.865 98.935 ;
		RECT	12.52 98.805 12.57 98.935 ;
		RECT	13.98 98.805 14.03 98.935 ;
		RECT	14.33 176.335 14.38 176.465 ;
		RECT	6.22 175.875 6.27 176.005 ;
		RECT	7.5 175.875 7.55 176.005 ;
		RECT	9.04 175.875 9.09 176.005 ;
		RECT	9.315 175.875 9.365 176.005 ;
		RECT	9.72 175.875 9.77 176.005 ;
		RECT	11.025 175.875 11.075 176.005 ;
		RECT	12.79 175.875 12.84 176.005 ;
		RECT	14.33 173.915 14.38 174.045 ;
		RECT	5.675 173.685 5.725 173.815 ;
		RECT	6.065 173.685 6.115 173.815 ;
		RECT	6.725 173.685 6.775 173.815 ;
		RECT	8.42 173.685 8.47 173.815 ;
		RECT	8.77 173.685 8.82 173.815 ;
		RECT	11.555 173.685 11.605 173.815 ;
		RECT	11.815 173.685 11.865 173.815 ;
		RECT	12.52 173.685 12.57 173.815 ;
		RECT	13.98 173.685 14.03 173.815 ;
		RECT	14.33 98.575 14.38 98.705 ;
		RECT	6.22 98.115 6.27 98.245 ;
		RECT	7.5 98.115 7.55 98.245 ;
		RECT	9.04 98.115 9.09 98.245 ;
		RECT	9.315 98.115 9.365 98.245 ;
		RECT	9.72 98.115 9.77 98.245 ;
		RECT	11.025 98.115 11.075 98.245 ;
		RECT	12.79 98.115 12.84 98.245 ;
		RECT	14.33 96.155 14.38 96.285 ;
		RECT	5.675 95.925 5.725 96.055 ;
		RECT	6.065 95.925 6.115 96.055 ;
		RECT	6.725 95.925 6.775 96.055 ;
		RECT	8.42 95.925 8.47 96.055 ;
		RECT	8.77 95.925 8.82 96.055 ;
		RECT	11.555 95.925 11.605 96.055 ;
		RECT	11.815 95.925 11.865 96.055 ;
		RECT	12.52 95.925 12.57 96.055 ;
		RECT	13.98 95.925 14.03 96.055 ;
		RECT	14.33 95.695 14.38 95.825 ;
		RECT	6.22 95.235 6.27 95.365 ;
		RECT	7.5 95.235 7.55 95.365 ;
		RECT	9.04 95.235 9.09 95.365 ;
		RECT	9.315 95.235 9.365 95.365 ;
		RECT	9.72 95.235 9.77 95.365 ;
		RECT	11.025 95.235 11.075 95.365 ;
		RECT	12.79 95.235 12.84 95.365 ;
		RECT	14.33 93.275 14.38 93.405 ;
		RECT	5.675 93.045 5.725 93.175 ;
		RECT	6.065 93.045 6.115 93.175 ;
		RECT	6.725 93.045 6.775 93.175 ;
		RECT	8.42 93.045 8.47 93.175 ;
		RECT	8.77 93.045 8.82 93.175 ;
		RECT	11.555 93.045 11.605 93.175 ;
		RECT	11.815 93.045 11.865 93.175 ;
		RECT	12.52 93.045 12.57 93.175 ;
		RECT	13.98 93.045 14.03 93.175 ;
		RECT	14.33 92.815 14.38 92.945 ;
		RECT	6.22 92.355 6.27 92.485 ;
		RECT	7.5 92.355 7.55 92.485 ;
		RECT	9.04 92.355 9.09 92.485 ;
		RECT	9.315 92.355 9.365 92.485 ;
		RECT	9.72 92.355 9.77 92.485 ;
		RECT	11.025 92.355 11.075 92.485 ;
		RECT	12.79 92.355 12.84 92.485 ;
		RECT	14.33 90.395 14.38 90.525 ;
		RECT	5.675 90.165 5.725 90.295 ;
		RECT	6.065 90.165 6.115 90.295 ;
		RECT	6.725 90.165 6.775 90.295 ;
		RECT	8.42 90.165 8.47 90.295 ;
		RECT	8.77 90.165 8.82 90.295 ;
		RECT	11.555 90.165 11.605 90.295 ;
		RECT	11.815 90.165 11.865 90.295 ;
		RECT	12.52 90.165 12.57 90.295 ;
		RECT	13.98 90.165 14.03 90.295 ;
		RECT	14.33 89.935 14.38 90.065 ;
		RECT	6.22 89.475 6.27 89.605 ;
		RECT	7.5 89.475 7.55 89.605 ;
		RECT	9.04 89.475 9.09 89.605 ;
		RECT	9.315 89.475 9.365 89.605 ;
		RECT	9.72 89.475 9.77 89.605 ;
		RECT	11.025 89.475 11.075 89.605 ;
		RECT	12.79 89.475 12.84 89.605 ;
		RECT	14.33 87.515 14.38 87.645 ;
		RECT	5.675 87.285 5.725 87.415 ;
		RECT	6.065 87.285 6.115 87.415 ;
		RECT	6.725 87.285 6.775 87.415 ;
		RECT	8.42 87.285 8.47 87.415 ;
		RECT	8.77 87.285 8.82 87.415 ;
		RECT	11.555 87.285 11.605 87.415 ;
		RECT	11.815 87.285 11.865 87.415 ;
		RECT	12.52 87.285 12.57 87.415 ;
		RECT	13.98 87.285 14.03 87.415 ;
		RECT	14.33 87.055 14.38 87.185 ;
		RECT	6.22 86.595 6.27 86.725 ;
		RECT	7.5 86.595 7.55 86.725 ;
		RECT	9.04 86.595 9.09 86.725 ;
		RECT	9.315 86.595 9.365 86.725 ;
		RECT	9.72 86.595 9.77 86.725 ;
		RECT	11.025 86.595 11.075 86.725 ;
		RECT	12.79 86.595 12.84 86.725 ;
		RECT	14.33 84.635 14.38 84.765 ;
		RECT	5.675 84.405 5.725 84.535 ;
		RECT	6.065 84.405 6.115 84.535 ;
		RECT	6.725 84.405 6.775 84.535 ;
		RECT	8.42 84.405 8.47 84.535 ;
		RECT	8.77 84.405 8.82 84.535 ;
		RECT	11.555 84.405 11.605 84.535 ;
		RECT	11.815 84.405 11.865 84.535 ;
		RECT	12.52 84.405 12.57 84.535 ;
		RECT	13.98 84.405 14.03 84.535 ;
		RECT	14.33 84.175 14.38 84.305 ;
		RECT	6.22 83.715 6.27 83.845 ;
		RECT	7.5 83.715 7.55 83.845 ;
		RECT	9.04 83.715 9.09 83.845 ;
		RECT	9.315 83.715 9.365 83.845 ;
		RECT	9.72 83.715 9.77 83.845 ;
		RECT	11.025 83.715 11.075 83.845 ;
		RECT	12.79 83.715 12.84 83.845 ;
		RECT	14.33 81.755 14.38 81.885 ;
		RECT	5.675 81.525 5.725 81.655 ;
		RECT	6.065 81.525 6.115 81.655 ;
		RECT	6.725 81.525 6.775 81.655 ;
		RECT	8.42 81.525 8.47 81.655 ;
		RECT	8.77 81.525 8.82 81.655 ;
		RECT	11.555 81.525 11.605 81.655 ;
		RECT	11.815 81.525 11.865 81.655 ;
		RECT	12.52 81.525 12.57 81.655 ;
		RECT	13.98 81.525 14.03 81.655 ;
		RECT	14.33 81.295 14.38 81.425 ;
		RECT	6.22 80.835 6.27 80.965 ;
		RECT	7.5 80.835 7.55 80.965 ;
		RECT	9.04 80.835 9.09 80.965 ;
		RECT	9.315 80.835 9.365 80.965 ;
		RECT	9.72 80.835 9.77 80.965 ;
		RECT	11.025 80.835 11.075 80.965 ;
		RECT	12.79 80.835 12.84 80.965 ;
		RECT	14.33 78.875 14.38 79.005 ;
		RECT	5.675 78.645 5.725 78.775 ;
		RECT	6.065 78.645 6.115 78.775 ;
		RECT	6.725 78.645 6.775 78.775 ;
		RECT	8.42 78.645 8.47 78.775 ;
		RECT	8.77 78.645 8.82 78.775 ;
		RECT	11.555 78.645 11.605 78.775 ;
		RECT	11.815 78.645 11.865 78.775 ;
		RECT	12.52 78.645 12.57 78.775 ;
		RECT	13.98 78.645 14.03 78.775 ;
		RECT	14.33 78.415 14.38 78.545 ;
		RECT	6.22 77.955 6.27 78.085 ;
		RECT	7.5 77.955 7.55 78.085 ;
		RECT	9.04 77.955 9.09 78.085 ;
		RECT	9.315 77.955 9.365 78.085 ;
		RECT	9.72 77.955 9.77 78.085 ;
		RECT	11.025 77.955 11.075 78.085 ;
		RECT	12.79 77.955 12.84 78.085 ;
		RECT	14.33 75.995 14.38 76.125 ;
		RECT	5.675 75.765 5.725 75.895 ;
		RECT	6.065 75.765 6.115 75.895 ;
		RECT	6.725 75.765 6.775 75.895 ;
		RECT	8.42 75.765 8.47 75.895 ;
		RECT	8.77 75.765 8.82 75.895 ;
		RECT	11.555 75.765 11.605 75.895 ;
		RECT	11.815 75.765 11.865 75.895 ;
		RECT	12.52 75.765 12.57 75.895 ;
		RECT	13.98 75.765 14.03 75.895 ;
		RECT	14.33 75.535 14.38 75.665 ;
		RECT	6.22 75.075 6.27 75.205 ;
		RECT	7.5 75.075 7.55 75.205 ;
		RECT	9.04 75.075 9.09 75.205 ;
		RECT	9.315 75.075 9.365 75.205 ;
		RECT	9.72 75.075 9.77 75.205 ;
		RECT	11.025 75.075 11.075 75.205 ;
		RECT	12.79 75.075 12.84 75.205 ;
		RECT	14.33 73.115 14.38 73.245 ;
		RECT	5.675 72.885 5.725 73.015 ;
		RECT	6.065 72.885 6.115 73.015 ;
		RECT	6.725 72.885 6.775 73.015 ;
		RECT	8.42 72.885 8.47 73.015 ;
		RECT	8.77 72.885 8.82 73.015 ;
		RECT	11.555 72.885 11.605 73.015 ;
		RECT	11.815 72.885 11.865 73.015 ;
		RECT	12.52 72.885 12.57 73.015 ;
		RECT	13.98 72.885 14.03 73.015 ;
		RECT	14.33 72.655 14.38 72.785 ;
		RECT	6.22 72.195 6.27 72.325 ;
		RECT	7.5 72.195 7.55 72.325 ;
		RECT	9.04 72.195 9.09 72.325 ;
		RECT	9.315 72.195 9.365 72.325 ;
		RECT	9.72 72.195 9.77 72.325 ;
		RECT	11.025 72.195 11.075 72.325 ;
		RECT	12.79 72.195 12.84 72.325 ;
		RECT	14.33 70.235 14.38 70.365 ;
		RECT	5.675 70.005 5.725 70.135 ;
		RECT	6.065 70.005 6.115 70.135 ;
		RECT	6.725 70.005 6.775 70.135 ;
		RECT	8.42 70.005 8.47 70.135 ;
		RECT	8.77 70.005 8.82 70.135 ;
		RECT	11.555 70.005 11.605 70.135 ;
		RECT	11.815 70.005 11.865 70.135 ;
		RECT	12.52 70.005 12.57 70.135 ;
		RECT	13.98 70.005 14.03 70.135 ;
		RECT	14.33 173.455 14.38 173.585 ;
		RECT	6.22 172.995 6.27 173.125 ;
		RECT	7.5 172.995 7.55 173.125 ;
		RECT	9.04 172.995 9.09 173.125 ;
		RECT	9.315 172.995 9.365 173.125 ;
		RECT	9.72 172.995 9.77 173.125 ;
		RECT	11.025 172.995 11.075 173.125 ;
		RECT	12.79 172.995 12.84 173.125 ;
		RECT	14.33 171.035 14.38 171.165 ;
		RECT	5.675 170.805 5.725 170.935 ;
		RECT	6.065 170.805 6.115 170.935 ;
		RECT	6.725 170.805 6.775 170.935 ;
		RECT	8.42 170.805 8.47 170.935 ;
		RECT	8.77 170.805 8.82 170.935 ;
		RECT	11.555 170.805 11.605 170.935 ;
		RECT	11.815 170.805 11.865 170.935 ;
		RECT	12.52 170.805 12.57 170.935 ;
		RECT	13.98 170.805 14.03 170.935 ;
		RECT	14.33 69.775 14.38 69.905 ;
		RECT	6.22 69.315 6.27 69.445 ;
		RECT	7.5 69.315 7.55 69.445 ;
		RECT	9.04 69.315 9.09 69.445 ;
		RECT	9.315 69.315 9.365 69.445 ;
		RECT	9.72 69.315 9.77 69.445 ;
		RECT	11.025 69.315 11.075 69.445 ;
		RECT	12.79 69.315 12.84 69.445 ;
		RECT	14.33 67.355 14.38 67.485 ;
		RECT	5.675 67.125 5.725 67.255 ;
		RECT	6.065 67.125 6.115 67.255 ;
		RECT	6.725 67.125 6.775 67.255 ;
		RECT	8.42 67.125 8.47 67.255 ;
		RECT	8.77 67.125 8.82 67.255 ;
		RECT	11.555 67.125 11.605 67.255 ;
		RECT	11.815 67.125 11.865 67.255 ;
		RECT	12.52 67.125 12.57 67.255 ;
		RECT	13.98 67.125 14.03 67.255 ;
		RECT	14.33 66.895 14.38 67.025 ;
		RECT	6.22 66.435 6.27 66.565 ;
		RECT	7.5 66.435 7.55 66.565 ;
		RECT	9.04 66.435 9.09 66.565 ;
		RECT	9.315 66.435 9.365 66.565 ;
		RECT	9.72 66.435 9.77 66.565 ;
		RECT	11.025 66.435 11.075 66.565 ;
		RECT	12.79 66.435 12.84 66.565 ;
		RECT	14.33 64.475 14.38 64.605 ;
		RECT	5.675 64.245 5.725 64.375 ;
		RECT	6.065 64.245 6.115 64.375 ;
		RECT	6.725 64.245 6.775 64.375 ;
		RECT	8.42 64.245 8.47 64.375 ;
		RECT	8.77 64.245 8.82 64.375 ;
		RECT	11.555 64.245 11.605 64.375 ;
		RECT	11.815 64.245 11.865 64.375 ;
		RECT	12.52 64.245 12.57 64.375 ;
		RECT	13.98 64.245 14.03 64.375 ;
		RECT	14.33 64.015 14.38 64.145 ;
		RECT	6.22 63.555 6.27 63.685 ;
		RECT	7.5 63.555 7.55 63.685 ;
		RECT	9.04 63.555 9.09 63.685 ;
		RECT	9.315 63.555 9.365 63.685 ;
		RECT	9.72 63.555 9.77 63.685 ;
		RECT	11.025 63.555 11.075 63.685 ;
		RECT	12.79 63.555 12.84 63.685 ;
		RECT	14.33 61.595 14.38 61.725 ;
		RECT	5.675 61.365 5.725 61.495 ;
		RECT	6.065 61.365 6.115 61.495 ;
		RECT	6.725 61.365 6.775 61.495 ;
		RECT	8.42 61.365 8.47 61.495 ;
		RECT	8.77 61.365 8.82 61.495 ;
		RECT	11.555 61.365 11.605 61.495 ;
		RECT	11.815 61.365 11.865 61.495 ;
		RECT	12.52 61.365 12.57 61.495 ;
		RECT	13.98 61.365 14.03 61.495 ;
		RECT	14.33 61.135 14.38 61.265 ;
		RECT	6.22 60.675 6.27 60.805 ;
		RECT	7.5 60.675 7.55 60.805 ;
		RECT	9.04 60.675 9.09 60.805 ;
		RECT	9.315 60.675 9.365 60.805 ;
		RECT	9.72 60.675 9.77 60.805 ;
		RECT	11.025 60.675 11.075 60.805 ;
		RECT	12.79 60.675 12.84 60.805 ;
		RECT	14.33 58.715 14.38 58.845 ;
		RECT	5.675 58.485 5.725 58.615 ;
		RECT	6.065 58.485 6.115 58.615 ;
		RECT	6.725 58.485 6.775 58.615 ;
		RECT	8.42 58.485 8.47 58.615 ;
		RECT	8.77 58.485 8.82 58.615 ;
		RECT	11.555 58.485 11.605 58.615 ;
		RECT	11.815 58.485 11.865 58.615 ;
		RECT	12.52 58.485 12.57 58.615 ;
		RECT	13.98 58.485 14.03 58.615 ;
		RECT	14.33 58.255 14.38 58.385 ;
		RECT	6.22 57.795 6.27 57.925 ;
		RECT	7.5 57.795 7.55 57.925 ;
		RECT	9.04 57.795 9.09 57.925 ;
		RECT	9.315 57.795 9.365 57.925 ;
		RECT	9.72 57.795 9.77 57.925 ;
		RECT	11.025 57.795 11.075 57.925 ;
		RECT	12.79 57.795 12.84 57.925 ;
		RECT	14.33 55.835 14.38 55.965 ;
		RECT	5.675 55.605 5.725 55.735 ;
		RECT	6.065 55.605 6.115 55.735 ;
		RECT	6.725 55.605 6.775 55.735 ;
		RECT	8.42 55.605 8.47 55.735 ;
		RECT	8.77 55.605 8.82 55.735 ;
		RECT	11.555 55.605 11.605 55.735 ;
		RECT	11.815 55.605 11.865 55.735 ;
		RECT	12.52 55.605 12.57 55.735 ;
		RECT	13.98 55.605 14.03 55.735 ;
		RECT	14.33 55.375 14.38 55.505 ;
		RECT	6.22 54.915 6.27 55.045 ;
		RECT	7.5 54.915 7.55 55.045 ;
		RECT	9.04 54.915 9.09 55.045 ;
		RECT	9.315 54.915 9.365 55.045 ;
		RECT	9.72 54.915 9.77 55.045 ;
		RECT	11.025 54.915 11.075 55.045 ;
		RECT	12.79 54.915 12.84 55.045 ;
		RECT	14.33 52.955 14.38 53.085 ;
		RECT	5.675 52.725 5.725 52.855 ;
		RECT	6.065 52.725 6.115 52.855 ;
		RECT	6.725 52.725 6.775 52.855 ;
		RECT	8.42 52.725 8.47 52.855 ;
		RECT	8.77 52.725 8.82 52.855 ;
		RECT	11.555 52.725 11.605 52.855 ;
		RECT	11.815 52.725 11.865 52.855 ;
		RECT	12.52 52.725 12.57 52.855 ;
		RECT	13.98 52.725 14.03 52.855 ;
		RECT	14.33 52.495 14.38 52.625 ;
		RECT	6.22 52.035 6.27 52.165 ;
		RECT	7.5 52.035 7.55 52.165 ;
		RECT	9.04 52.035 9.09 52.165 ;
		RECT	9.315 52.035 9.365 52.165 ;
		RECT	9.72 52.035 9.77 52.165 ;
		RECT	11.025 52.035 11.075 52.165 ;
		RECT	12.79 52.035 12.84 52.165 ;
		RECT	14.33 50.075 14.38 50.205 ;
		RECT	5.675 49.845 5.725 49.975 ;
		RECT	6.065 49.845 6.115 49.975 ;
		RECT	6.725 49.845 6.775 49.975 ;
		RECT	8.42 49.845 8.47 49.975 ;
		RECT	8.77 49.845 8.82 49.975 ;
		RECT	11.555 49.845 11.605 49.975 ;
		RECT	11.815 49.845 11.865 49.975 ;
		RECT	12.52 49.845 12.57 49.975 ;
		RECT	13.98 49.845 14.03 49.975 ;
		RECT	14.33 49.615 14.38 49.745 ;
		RECT	6.22 49.155 6.27 49.285 ;
		RECT	7.5 49.155 7.55 49.285 ;
		RECT	9.04 49.155 9.09 49.285 ;
		RECT	9.315 49.155 9.365 49.285 ;
		RECT	9.72 49.155 9.77 49.285 ;
		RECT	11.025 49.155 11.075 49.285 ;
		RECT	12.79 49.155 12.84 49.285 ;
		RECT	14.33 47.195 14.38 47.325 ;
		RECT	5.675 46.965 5.725 47.095 ;
		RECT	6.065 46.965 6.115 47.095 ;
		RECT	6.725 46.965 6.775 47.095 ;
		RECT	8.42 46.965 8.47 47.095 ;
		RECT	8.77 46.965 8.82 47.095 ;
		RECT	11.555 46.965 11.605 47.095 ;
		RECT	11.815 46.965 11.865 47.095 ;
		RECT	12.52 46.965 12.57 47.095 ;
		RECT	13.98 46.965 14.03 47.095 ;
		RECT	14.33 46.735 14.38 46.865 ;
		RECT	6.22 46.275 6.27 46.405 ;
		RECT	7.5 46.275 7.55 46.405 ;
		RECT	9.04 46.275 9.09 46.405 ;
		RECT	9.315 46.275 9.365 46.405 ;
		RECT	9.72 46.275 9.77 46.405 ;
		RECT	11.025 46.275 11.075 46.405 ;
		RECT	12.79 46.275 12.84 46.405 ;
		RECT	14.33 44.315 14.38 44.445 ;
		RECT	5.675 44.085 5.725 44.215 ;
		RECT	6.065 44.085 6.115 44.215 ;
		RECT	6.725 44.085 6.775 44.215 ;
		RECT	8.42 44.085 8.47 44.215 ;
		RECT	8.77 44.085 8.82 44.215 ;
		RECT	11.555 44.085 11.605 44.215 ;
		RECT	11.815 44.085 11.865 44.215 ;
		RECT	12.52 44.085 12.57 44.215 ;
		RECT	13.98 44.085 14.03 44.215 ;
		RECT	14.33 43.855 14.38 43.985 ;
		RECT	6.22 43.395 6.27 43.525 ;
		RECT	7.5 43.395 7.55 43.525 ;
		RECT	9.04 43.395 9.09 43.525 ;
		RECT	9.315 43.395 9.365 43.525 ;
		RECT	9.72 43.395 9.77 43.525 ;
		RECT	11.025 43.395 11.075 43.525 ;
		RECT	12.79 43.395 12.84 43.525 ;
		RECT	14.33 41.435 14.38 41.565 ;
		RECT	5.675 41.205 5.725 41.335 ;
		RECT	6.065 41.205 6.115 41.335 ;
		RECT	6.725 41.205 6.775 41.335 ;
		RECT	8.42 41.205 8.47 41.335 ;
		RECT	8.77 41.205 8.82 41.335 ;
		RECT	11.555 41.205 11.605 41.335 ;
		RECT	11.815 41.205 11.865 41.335 ;
		RECT	12.52 41.205 12.57 41.335 ;
		RECT	13.98 41.205 14.03 41.335 ;
		RECT	14.33 170.575 14.38 170.705 ;
		RECT	6.22 170.115 6.27 170.245 ;
		RECT	7.5 170.115 7.55 170.245 ;
		RECT	9.04 170.115 9.09 170.245 ;
		RECT	9.315 170.115 9.365 170.245 ;
		RECT	9.72 170.115 9.77 170.245 ;
		RECT	11.025 170.115 11.075 170.245 ;
		RECT	12.79 170.115 12.84 170.245 ;
		RECT	14.33 168.155 14.38 168.285 ;
		RECT	5.675 167.925 5.725 168.055 ;
		RECT	6.065 167.925 6.115 168.055 ;
		RECT	6.725 167.925 6.775 168.055 ;
		RECT	8.42 167.925 8.47 168.055 ;
		RECT	8.77 167.925 8.82 168.055 ;
		RECT	11.555 167.925 11.605 168.055 ;
		RECT	11.815 167.925 11.865 168.055 ;
		RECT	12.52 167.925 12.57 168.055 ;
		RECT	13.98 167.925 14.03 168.055 ;
		RECT	14.33 40.975 14.38 41.105 ;
		RECT	6.22 40.515 6.27 40.645 ;
		RECT	7.5 40.515 7.55 40.645 ;
		RECT	9.04 40.515 9.09 40.645 ;
		RECT	9.315 40.515 9.365 40.645 ;
		RECT	9.72 40.515 9.77 40.645 ;
		RECT	11.025 40.515 11.075 40.645 ;
		RECT	12.79 40.515 12.84 40.645 ;
		RECT	14.33 38.555 14.38 38.685 ;
		RECT	5.675 38.325 5.725 38.455 ;
		RECT	6.065 38.325 6.115 38.455 ;
		RECT	6.725 38.325 6.775 38.455 ;
		RECT	8.42 38.325 8.47 38.455 ;
		RECT	8.77 38.325 8.82 38.455 ;
		RECT	11.555 38.325 11.605 38.455 ;
		RECT	11.815 38.325 11.865 38.455 ;
		RECT	12.52 38.325 12.57 38.455 ;
		RECT	13.98 38.325 14.03 38.455 ;
		RECT	14.33 38.095 14.38 38.225 ;
		RECT	6.22 37.635 6.27 37.765 ;
		RECT	7.5 37.635 7.55 37.765 ;
		RECT	9.04 37.635 9.09 37.765 ;
		RECT	9.315 37.635 9.365 37.765 ;
		RECT	9.72 37.635 9.77 37.765 ;
		RECT	11.025 37.635 11.075 37.765 ;
		RECT	12.79 37.635 12.84 37.765 ;
		RECT	14.33 35.675 14.38 35.805 ;
		RECT	5.675 35.445 5.725 35.575 ;
		RECT	6.065 35.445 6.115 35.575 ;
		RECT	6.725 35.445 6.775 35.575 ;
		RECT	8.42 35.445 8.47 35.575 ;
		RECT	8.77 35.445 8.82 35.575 ;
		RECT	11.555 35.445 11.605 35.575 ;
		RECT	11.815 35.445 11.865 35.575 ;
		RECT	12.52 35.445 12.57 35.575 ;
		RECT	13.98 35.445 14.03 35.575 ;
		RECT	14.33 35.215 14.38 35.345 ;
		RECT	6.22 34.755 6.27 34.885 ;
		RECT	7.5 34.755 7.55 34.885 ;
		RECT	9.04 34.755 9.09 34.885 ;
		RECT	9.315 34.755 9.365 34.885 ;
		RECT	9.72 34.755 9.77 34.885 ;
		RECT	11.025 34.755 11.075 34.885 ;
		RECT	12.79 34.755 12.84 34.885 ;
		RECT	14.33 32.795 14.38 32.925 ;
		RECT	5.675 32.565 5.725 32.695 ;
		RECT	6.065 32.565 6.115 32.695 ;
		RECT	6.725 32.565 6.775 32.695 ;
		RECT	8.42 32.565 8.47 32.695 ;
		RECT	8.77 32.565 8.82 32.695 ;
		RECT	11.555 32.565 11.605 32.695 ;
		RECT	11.815 32.565 11.865 32.695 ;
		RECT	12.52 32.565 12.57 32.695 ;
		RECT	13.98 32.565 14.03 32.695 ;
		RECT	14.33 32.335 14.38 32.465 ;
		RECT	6.22 31.875 6.27 32.005 ;
		RECT	7.5 31.875 7.55 32.005 ;
		RECT	9.04 31.875 9.09 32.005 ;
		RECT	9.315 31.875 9.365 32.005 ;
		RECT	9.72 31.875 9.77 32.005 ;
		RECT	11.025 31.875 11.075 32.005 ;
		RECT	12.79 31.875 12.84 32.005 ;
		RECT	14.33 29.915 14.38 30.045 ;
		RECT	5.675 29.685 5.725 29.815 ;
		RECT	6.065 29.685 6.115 29.815 ;
		RECT	6.725 29.685 6.775 29.815 ;
		RECT	8.42 29.685 8.47 29.815 ;
		RECT	8.77 29.685 8.82 29.815 ;
		RECT	11.555 29.685 11.605 29.815 ;
		RECT	11.815 29.685 11.865 29.815 ;
		RECT	12.52 29.685 12.57 29.815 ;
		RECT	13.98 29.685 14.03 29.815 ;
		RECT	14.33 29.455 14.38 29.585 ;
		RECT	6.22 28.995 6.27 29.125 ;
		RECT	7.5 28.995 7.55 29.125 ;
		RECT	9.04 28.995 9.09 29.125 ;
		RECT	9.315 28.995 9.365 29.125 ;
		RECT	9.72 28.995 9.77 29.125 ;
		RECT	11.025 28.995 11.075 29.125 ;
		RECT	12.79 28.995 12.84 29.125 ;
		RECT	14.33 27.035 14.38 27.165 ;
		RECT	5.675 26.805 5.725 26.935 ;
		RECT	6.065 26.805 6.115 26.935 ;
		RECT	6.725 26.805 6.775 26.935 ;
		RECT	8.42 26.805 8.47 26.935 ;
		RECT	8.77 26.805 8.82 26.935 ;
		RECT	11.555 26.805 11.605 26.935 ;
		RECT	11.815 26.805 11.865 26.935 ;
		RECT	12.52 26.805 12.57 26.935 ;
		RECT	13.98 26.805 14.03 26.935 ;
		RECT	14.33 26.575 14.38 26.705 ;
		RECT	6.22 26.115 6.27 26.245 ;
		RECT	7.5 26.115 7.55 26.245 ;
		RECT	9.04 26.115 9.09 26.245 ;
		RECT	9.315 26.115 9.365 26.245 ;
		RECT	9.72 26.115 9.77 26.245 ;
		RECT	11.025 26.115 11.075 26.245 ;
		RECT	12.79 26.115 12.84 26.245 ;
		RECT	14.33 24.155 14.38 24.285 ;
		RECT	5.675 23.925 5.725 24.055 ;
		RECT	6.065 23.925 6.115 24.055 ;
		RECT	6.725 23.925 6.775 24.055 ;
		RECT	8.42 23.925 8.47 24.055 ;
		RECT	8.77 23.925 8.82 24.055 ;
		RECT	11.555 23.925 11.605 24.055 ;
		RECT	11.815 23.925 11.865 24.055 ;
		RECT	12.52 23.925 12.57 24.055 ;
		RECT	13.98 23.925 14.03 24.055 ;
		RECT	14.33 23.695 14.38 23.825 ;
		RECT	6.22 23.235 6.27 23.365 ;
		RECT	7.5 23.235 7.55 23.365 ;
		RECT	9.04 23.235 9.09 23.365 ;
		RECT	9.315 23.235 9.365 23.365 ;
		RECT	9.72 23.235 9.77 23.365 ;
		RECT	11.025 23.235 11.075 23.365 ;
		RECT	12.79 23.235 12.84 23.365 ;
		RECT	14.33 21.275 14.38 21.405 ;
		RECT	5.675 21.045 5.725 21.175 ;
		RECT	6.065 21.045 6.115 21.175 ;
		RECT	6.725 21.045 6.775 21.175 ;
		RECT	8.42 21.045 8.47 21.175 ;
		RECT	8.77 21.045 8.82 21.175 ;
		RECT	11.555 21.045 11.605 21.175 ;
		RECT	11.815 21.045 11.865 21.175 ;
		RECT	12.52 21.045 12.57 21.175 ;
		RECT	13.98 21.045 14.03 21.175 ;
		RECT	14.33 20.815 14.38 20.945 ;
		RECT	6.22 20.355 6.27 20.485 ;
		RECT	7.5 20.355 7.55 20.485 ;
		RECT	9.04 20.355 9.09 20.485 ;
		RECT	9.315 20.355 9.365 20.485 ;
		RECT	9.72 20.355 9.77 20.485 ;
		RECT	11.025 20.355 11.075 20.485 ;
		RECT	12.79 20.355 12.84 20.485 ;
		RECT	14.33 18.395 14.38 18.525 ;
		RECT	5.675 18.165 5.725 18.295 ;
		RECT	6.065 18.165 6.115 18.295 ;
		RECT	6.725 18.165 6.775 18.295 ;
		RECT	8.42 18.165 8.47 18.295 ;
		RECT	8.77 18.165 8.82 18.295 ;
		RECT	11.555 18.165 11.605 18.295 ;
		RECT	11.815 18.165 11.865 18.295 ;
		RECT	12.52 18.165 12.57 18.295 ;
		RECT	13.98 18.165 14.03 18.295 ;
		RECT	14.33 17.935 14.38 18.065 ;
		RECT	6.22 17.475 6.27 17.605 ;
		RECT	7.5 17.475 7.55 17.605 ;
		RECT	9.04 17.475 9.09 17.605 ;
		RECT	9.315 17.475 9.365 17.605 ;
		RECT	9.72 17.475 9.77 17.605 ;
		RECT	11.025 17.475 11.075 17.605 ;
		RECT	12.79 17.475 12.84 17.605 ;
		RECT	14.33 15.515 14.38 15.645 ;
		RECT	5.675 15.285 5.725 15.415 ;
		RECT	6.065 15.285 6.115 15.415 ;
		RECT	6.725 15.285 6.775 15.415 ;
		RECT	8.42 15.285 8.47 15.415 ;
		RECT	8.77 15.285 8.82 15.415 ;
		RECT	11.555 15.285 11.605 15.415 ;
		RECT	11.815 15.285 11.865 15.415 ;
		RECT	12.52 15.285 12.57 15.415 ;
		RECT	13.98 15.285 14.03 15.415 ;
		RECT	14.33 15.055 14.38 15.185 ;
		RECT	6.22 14.595 6.27 14.725 ;
		RECT	7.5 14.595 7.55 14.725 ;
		RECT	9.04 14.595 9.09 14.725 ;
		RECT	9.315 14.595 9.365 14.725 ;
		RECT	9.72 14.595 9.77 14.725 ;
		RECT	11.025 14.595 11.075 14.725 ;
		RECT	12.79 14.595 12.84 14.725 ;
		RECT	14.33 12.635 14.38 12.765 ;
		RECT	5.675 12.405 5.725 12.535 ;
		RECT	6.065 12.405 6.115 12.535 ;
		RECT	6.725 12.405 6.775 12.535 ;
		RECT	8.42 12.405 8.47 12.535 ;
		RECT	8.77 12.405 8.82 12.535 ;
		RECT	11.555 12.405 11.605 12.535 ;
		RECT	11.815 12.405 11.865 12.535 ;
		RECT	12.52 12.405 12.57 12.535 ;
		RECT	13.98 12.405 14.03 12.535 ;
		RECT	14.33 167.695 14.38 167.825 ;
		RECT	6.22 167.235 6.27 167.365 ;
		RECT	7.5 167.235 7.55 167.365 ;
		RECT	9.04 167.235 9.09 167.365 ;
		RECT	9.315 167.235 9.365 167.365 ;
		RECT	9.72 167.235 9.77 167.365 ;
		RECT	11.025 167.235 11.075 167.365 ;
		RECT	12.79 167.235 12.84 167.365 ;
		RECT	14.33 165.275 14.38 165.405 ;
		RECT	5.675 165.045 5.725 165.175 ;
		RECT	6.065 165.045 6.115 165.175 ;
		RECT	6.725 165.045 6.775 165.175 ;
		RECT	8.42 165.045 8.47 165.175 ;
		RECT	8.77 165.045 8.82 165.175 ;
		RECT	11.555 165.045 11.605 165.175 ;
		RECT	11.815 165.045 11.865 165.175 ;
		RECT	12.52 165.045 12.57 165.175 ;
		RECT	13.98 165.045 14.03 165.175 ;
		RECT	14.33 12.175 14.38 12.305 ;
		RECT	6.22 11.715 6.27 11.845 ;
		RECT	7.5 11.715 7.55 11.845 ;
		RECT	9.04 11.715 9.09 11.845 ;
		RECT	9.315 11.715 9.365 11.845 ;
		RECT	9.72 11.715 9.77 11.845 ;
		RECT	11.025 11.715 11.075 11.845 ;
		RECT	12.79 11.715 12.84 11.845 ;
		RECT	14.33 9.755 14.38 9.885 ;
		RECT	5.675 9.525 5.725 9.655 ;
		RECT	6.065 9.525 6.115 9.655 ;
		RECT	6.725 9.525 6.775 9.655 ;
		RECT	8.42 9.525 8.47 9.655 ;
		RECT	8.77 9.525 8.82 9.655 ;
		RECT	11.555 9.525 11.605 9.655 ;
		RECT	11.815 9.525 11.865 9.655 ;
		RECT	12.52 9.525 12.57 9.655 ;
		RECT	13.98 9.525 14.03 9.655 ;
		RECT	14.33 9.295 14.38 9.425 ;
		RECT	6.22 8.835 6.27 8.965 ;
		RECT	7.5 8.835 7.55 8.965 ;
		RECT	9.04 8.835 9.09 8.965 ;
		RECT	9.315 8.835 9.365 8.965 ;
		RECT	9.72 8.835 9.77 8.965 ;
		RECT	11.025 8.835 11.075 8.965 ;
		RECT	12.79 8.835 12.84 8.965 ;
		RECT	14.33 6.875 14.38 7.005 ;
		RECT	5.675 6.645 5.725 6.775 ;
		RECT	6.065 6.645 6.115 6.775 ;
		RECT	6.725 6.645 6.775 6.775 ;
		RECT	8.42 6.645 8.47 6.775 ;
		RECT	8.77 6.645 8.82 6.775 ;
		RECT	11.555 6.645 11.605 6.775 ;
		RECT	11.815 6.645 11.865 6.775 ;
		RECT	12.52 6.645 12.57 6.775 ;
		RECT	13.98 6.645 14.03 6.775 ;
		RECT	14.33 6.415 14.38 6.545 ;
		RECT	6.22 5.955 6.27 6.085 ;
		RECT	7.5 5.955 7.55 6.085 ;
		RECT	9.04 5.955 9.09 6.085 ;
		RECT	9.315 5.955 9.365 6.085 ;
		RECT	9.72 5.955 9.77 6.085 ;
		RECT	11.025 5.955 11.075 6.085 ;
		RECT	12.79 5.955 12.84 6.085 ;
		RECT	14.33 3.995 14.38 4.125 ;
		RECT	5.675 3.765 5.725 3.895 ;
		RECT	6.065 3.765 6.115 3.895 ;
		RECT	6.725 3.765 6.775 3.895 ;
		RECT	8.42 3.765 8.47 3.895 ;
		RECT	8.77 3.765 8.82 3.895 ;
		RECT	11.555 3.765 11.605 3.895 ;
		RECT	11.815 3.765 11.865 3.895 ;
		RECT	12.52 3.765 12.57 3.895 ;
		RECT	13.98 3.765 14.03 3.895 ;
		RECT	14.33 164.815 14.38 164.945 ;
		RECT	6.22 164.355 6.27 164.485 ;
		RECT	7.5 164.355 7.55 164.485 ;
		RECT	9.04 164.355 9.09 164.485 ;
		RECT	9.315 164.355 9.365 164.485 ;
		RECT	9.72 164.355 9.77 164.485 ;
		RECT	11.025 164.355 11.075 164.485 ;
		RECT	12.79 164.355 12.84 164.485 ;
		RECT	14.33 162.395 14.38 162.525 ;
		RECT	5.675 162.165 5.725 162.295 ;
		RECT	6.065 162.165 6.115 162.295 ;
		RECT	6.725 162.165 6.775 162.295 ;
		RECT	8.42 162.165 8.47 162.295 ;
		RECT	8.77 162.165 8.82 162.295 ;
		RECT	11.555 162.165 11.605 162.295 ;
		RECT	11.815 162.165 11.865 162.295 ;
		RECT	12.52 162.165 12.57 162.295 ;
		RECT	13.98 162.165 14.03 162.295 ;
		RECT	14.33 161.935 14.38 162.065 ;
		RECT	6.22 161.475 6.27 161.605 ;
		RECT	7.5 161.475 7.55 161.605 ;
		RECT	9.04 161.475 9.09 161.605 ;
		RECT	9.315 161.475 9.365 161.605 ;
		RECT	9.72 161.475 9.77 161.605 ;
		RECT	11.025 161.475 11.075 161.605 ;
		RECT	12.79 161.475 12.84 161.605 ;
		RECT	14.33 159.515 14.38 159.645 ;
		RECT	5.675 159.285 5.725 159.415 ;
		RECT	6.065 159.285 6.115 159.415 ;
		RECT	6.725 159.285 6.775 159.415 ;
		RECT	8.42 159.285 8.47 159.415 ;
		RECT	8.77 159.285 8.82 159.415 ;
		RECT	11.555 159.285 11.605 159.415 ;
		RECT	11.815 159.285 11.865 159.415 ;
		RECT	12.52 159.285 12.57 159.415 ;
		RECT	13.98 159.285 14.03 159.415 ;
		RECT	14.33 159.055 14.38 159.185 ;
		RECT	6.22 158.595 6.27 158.725 ;
		RECT	7.5 158.595 7.55 158.725 ;
		RECT	9.04 158.595 9.09 158.725 ;
		RECT	9.315 158.595 9.365 158.725 ;
		RECT	9.72 158.595 9.77 158.725 ;
		RECT	11.025 158.595 11.075 158.725 ;
		RECT	12.79 158.595 12.84 158.725 ;
		RECT	14.33 156.635 14.38 156.765 ;
		RECT	5.675 156.405 5.725 156.535 ;
		RECT	6.065 156.405 6.115 156.535 ;
		RECT	6.725 156.405 6.775 156.535 ;
		RECT	8.42 156.405 8.47 156.535 ;
		RECT	8.77 156.405 8.82 156.535 ;
		RECT	11.555 156.405 11.605 156.535 ;
		RECT	11.815 156.405 11.865 156.535 ;
		RECT	12.52 156.405 12.57 156.535 ;
		RECT	13.98 156.405 14.03 156.535 ;
		RECT	14.33 3.535 14.38 3.665 ;
		RECT	6.22 3.075 6.27 3.205 ;
		RECT	7.5 3.075 7.55 3.205 ;
		RECT	9.04 3.075 9.09 3.205 ;
		RECT	9.315 3.075 9.365 3.205 ;
		RECT	9.72 3.075 9.77 3.205 ;
		RECT	11.025 3.075 11.075 3.205 ;
		RECT	12.79 3.075 12.84 3.205 ;
		RECT	14.33 1.115 14.38 1.245 ;
		RECT	5.675 0.885 5.725 1.015 ;
		RECT	6.065 0.885 6.115 1.015 ;
		RECT	6.725 0.885 6.775 1.015 ;
		RECT	8.42 0.885 8.47 1.015 ;
		RECT	8.77 0.885 8.82 1.015 ;
		RECT	11.555 0.885 11.605 1.015 ;
		RECT	11.815 0.885 11.865 1.015 ;
		RECT	12.52 0.885 12.57 1.015 ;
		RECT	13.98 0.885 14.03 1.015 ;
		RECT	14.33 184.975 14.38 185.105 ;
		RECT	6.22 184.515 6.27 184.645 ;
		RECT	7.5 184.515 7.55 184.645 ;
		RECT	9.04 184.515 9.09 184.645 ;
		RECT	9.315 184.515 9.365 184.645 ;
		RECT	9.72 184.515 9.77 184.645 ;
		RECT	11.025 184.515 11.075 184.645 ;
		RECT	12.79 184.515 12.84 184.645 ;
		RECT	14.33 182.555 14.38 182.685 ;
		RECT	5.675 182.325 5.725 182.455 ;
		RECT	6.065 182.325 6.115 182.455 ;
		RECT	6.725 182.325 6.775 182.455 ;
		RECT	8.42 182.325 8.47 182.455 ;
		RECT	8.77 182.325 8.82 182.455 ;
		RECT	11.555 182.325 11.605 182.455 ;
		RECT	11.815 182.325 11.865 182.455 ;
		RECT	12.52 182.325 12.57 182.455 ;
		RECT	13.98 182.325 14.03 182.455 ;
		RECT	13.98 0.195 14.03 0.325 ;
		RECT	3.06 0.655 3.11 0.785 ;
		RECT	1.57 0.195 1.62 0.325 ;
		RECT	2.485 0.195 2.665 0.325 ;
		RECT	3.84 0.195 3.89 0.325 ;
		RECT	7.19 0.195 7.24 0.325 ;
		RECT	14.14 0.195 14.19 0.325 ;
		RECT	13.8 0.425 13.85 0.555 ;
		RECT	8.56 0.655 8.61 0.785 ;
		RECT	10.27 0.655 10.32 0.785 ;
		RECT	0.435 0.655 0.485 0.785 ;
		RECT	0.62 0.195 0.67 0.325 ;
		RECT	3.65 0.195 3.7 0.325 ;
		RECT	2.18 0.655 2.23 0.785 ;
		RECT	0.9 179.445 0.95 179.575 ;
		RECT	0.9 153.525 0.95 153.655 ;
		RECT	0.9 150.645 0.95 150.775 ;
		RECT	0.9 147.765 0.95 147.895 ;
		RECT	0.9 144.885 0.95 145.015 ;
		RECT	0.9 142.005 0.95 142.135 ;
		RECT	0.9 139.125 0.95 139.255 ;
		RECT	0.9 136.245 0.95 136.375 ;
		RECT	0.9 133.365 0.95 133.495 ;
		RECT	0.9 130.485 0.95 130.615 ;
		RECT	0.9 127.605 0.95 127.735 ;
		RECT	0.9 176.565 0.95 176.695 ;
		RECT	0.9 124.725 0.95 124.855 ;
		RECT	0.9 121.845 0.95 121.975 ;
		RECT	0.9 118.965 0.95 119.095 ;
		RECT	0.9 116.085 0.95 116.215 ;
		RECT	0.9 113.205 0.95 113.335 ;
		RECT	0.9 110.325 0.95 110.455 ;
		RECT	0.9 107.445 0.95 107.575 ;
		RECT	0.9 104.565 0.95 104.695 ;
		RECT	0.9 101.685 0.95 101.815 ;
		RECT	0.9 98.805 0.95 98.935 ;
		RECT	0.9 173.685 0.95 173.815 ;
		RECT	0.9 95.925 0.95 96.055 ;
		RECT	0.9 93.045 0.95 93.175 ;
		RECT	0.9 90.165 0.95 90.295 ;
		RECT	0.9 87.285 0.95 87.415 ;
		RECT	0.9 84.405 0.95 84.535 ;
		RECT	0.9 81.525 0.95 81.655 ;
		RECT	0.9 78.645 0.95 78.775 ;
		RECT	0.9 75.765 0.95 75.895 ;
		RECT	0.9 72.885 0.95 73.015 ;
		RECT	0.9 70.005 0.95 70.135 ;
		RECT	0.9 170.805 0.95 170.935 ;
		RECT	0.9 67.125 0.95 67.255 ;
		RECT	0.9 64.245 0.95 64.375 ;
		RECT	0.9 61.365 0.95 61.495 ;
		RECT	0.9 58.485 0.95 58.615 ;
		RECT	0.9 55.605 0.95 55.735 ;
		RECT	0.9 52.725 0.95 52.855 ;
		RECT	0.9 49.845 0.95 49.975 ;
		RECT	0.9 46.965 0.95 47.095 ;
		RECT	0.9 44.085 0.95 44.215 ;
		RECT	0.9 41.205 0.95 41.335 ;
		RECT	0.9 167.925 0.95 168.055 ;
		RECT	0.9 38.325 0.95 38.455 ;
		RECT	0.9 35.445 0.95 35.575 ;
		RECT	0.9 32.565 0.95 32.695 ;
		RECT	0.9 29.685 0.95 29.815 ;
		RECT	0.9 26.805 0.95 26.935 ;
		RECT	0.9 23.925 0.95 24.055 ;
		RECT	0.9 21.045 0.95 21.175 ;
		RECT	0.9 18.165 0.95 18.295 ;
		RECT	0.9 15.285 0.95 15.415 ;
		RECT	0.9 12.405 0.95 12.535 ;
		RECT	0.9 165.045 0.95 165.175 ;
		RECT	0.9 9.525 0.95 9.655 ;
		RECT	0.9 6.645 0.95 6.775 ;
		RECT	0.9 3.765 0.95 3.895 ;
		RECT	0.9 162.165 0.95 162.295 ;
		RECT	0.9 159.285 0.95 159.415 ;
		RECT	0.9 156.405 0.95 156.535 ;
		RECT	0.9 0.885 0.95 1.015 ;
		RECT	0.9 182.325 0.95 182.455 ;
		RECT	2.18 184.975 2.23 185.105 ;
		RECT	2.18 182.555 2.23 182.685 ;
		RECT	2.18 156.175 2.23 156.305 ;
		RECT	2.18 153.755 2.23 153.885 ;
		RECT	2.18 153.295 2.23 153.425 ;
		RECT	2.18 150.875 2.23 151.005 ;
		RECT	2.18 150.415 2.23 150.545 ;
		RECT	2.18 147.995 2.23 148.125 ;
		RECT	2.18 147.535 2.23 147.665 ;
		RECT	2.18 145.115 2.23 145.245 ;
		RECT	2.18 144.655 2.23 144.785 ;
		RECT	2.18 142.235 2.23 142.365 ;
		RECT	2.18 141.775 2.23 141.905 ;
		RECT	2.18 139.355 2.23 139.485 ;
		RECT	2.18 138.895 2.23 139.025 ;
		RECT	2.18 136.475 2.23 136.605 ;
		RECT	2.18 136.015 2.23 136.145 ;
		RECT	2.18 133.595 2.23 133.725 ;
		RECT	2.18 133.135 2.23 133.265 ;
		RECT	2.18 130.715 2.23 130.845 ;
		RECT	2.18 130.255 2.23 130.385 ;
		RECT	2.18 127.835 2.23 127.965 ;
		RECT	2.18 182.095 2.23 182.225 ;
		RECT	2.18 179.675 2.23 179.805 ;
		RECT	2.18 127.375 2.23 127.505 ;
		RECT	2.18 124.955 2.23 125.085 ;
		RECT	2.18 124.495 2.23 124.625 ;
		RECT	2.18 122.075 2.23 122.205 ;
		RECT	2.18 121.615 2.23 121.745 ;
		RECT	2.18 119.195 2.23 119.325 ;
		RECT	2.18 118.735 2.23 118.865 ;
		RECT	2.18 116.315 2.23 116.445 ;
		RECT	2.18 115.855 2.23 115.985 ;
		RECT	2.18 113.435 2.23 113.565 ;
		RECT	2.18 112.975 2.23 113.105 ;
		RECT	2.18 110.555 2.23 110.685 ;
		RECT	2.18 110.095 2.23 110.225 ;
		RECT	2.18 107.675 2.23 107.805 ;
		RECT	2.18 107.215 2.23 107.345 ;
		RECT	2.18 104.795 2.23 104.925 ;
		RECT	2.18 104.335 2.23 104.465 ;
		RECT	2.18 101.915 2.23 102.045 ;
		RECT	2.18 101.455 2.23 101.585 ;
		RECT	2.18 99.035 2.23 99.165 ;
		RECT	2.18 179.215 2.23 179.345 ;
		RECT	2.18 176.795 2.23 176.925 ;
		RECT	2.18 98.575 2.23 98.705 ;
		RECT	2.18 96.155 2.23 96.285 ;
		RECT	2.18 95.695 2.23 95.825 ;
		RECT	2.18 93.275 2.23 93.405 ;
		RECT	2.18 92.815 2.23 92.945 ;
		RECT	2.18 90.395 2.23 90.525 ;
		RECT	2.18 89.935 2.23 90.065 ;
		RECT	2.18 87.515 2.23 87.645 ;
		RECT	2.18 87.055 2.23 87.185 ;
		RECT	2.18 84.635 2.23 84.765 ;
		RECT	2.18 84.175 2.23 84.305 ;
		RECT	2.18 81.755 2.23 81.885 ;
		RECT	2.18 81.295 2.23 81.425 ;
		RECT	2.18 78.875 2.23 79.005 ;
		RECT	2.18 78.415 2.23 78.545 ;
		RECT	2.18 75.995 2.23 76.125 ;
		RECT	2.18 75.535 2.23 75.665 ;
		RECT	2.18 73.115 2.23 73.245 ;
		RECT	2.18 72.655 2.23 72.785 ;
		RECT	2.18 70.235 2.23 70.365 ;
		RECT	2.18 176.335 2.23 176.465 ;
		RECT	2.18 173.915 2.23 174.045 ;
		RECT	2.18 69.775 2.23 69.905 ;
		RECT	2.18 67.355 2.23 67.485 ;
		RECT	2.18 66.895 2.23 67.025 ;
		RECT	2.18 64.475 2.23 64.605 ;
		RECT	2.18 64.015 2.23 64.145 ;
		RECT	2.18 61.595 2.23 61.725 ;
		RECT	2.18 61.135 2.23 61.265 ;
		RECT	2.18 58.715 2.23 58.845 ;
		RECT	2.18 58.255 2.23 58.385 ;
		RECT	2.18 55.835 2.23 55.965 ;
		RECT	2.18 55.375 2.23 55.505 ;
		RECT	2.18 52.955 2.23 53.085 ;
		RECT	2.18 52.495 2.23 52.625 ;
		RECT	2.18 50.075 2.23 50.205 ;
		RECT	2.18 49.615 2.23 49.745 ;
		RECT	2.18 47.195 2.23 47.325 ;
		RECT	2.18 46.735 2.23 46.865 ;
		RECT	2.18 44.315 2.23 44.445 ;
		RECT	2.18 43.855 2.23 43.985 ;
		RECT	2.18 41.435 2.23 41.565 ;
		RECT	2.18 173.455 2.23 173.585 ;
		RECT	2.18 171.035 2.23 171.165 ;
		RECT	2.18 40.975 2.23 41.105 ;
		RECT	2.18 38.555 2.23 38.685 ;
		RECT	2.18 38.095 2.23 38.225 ;
		RECT	2.18 35.675 2.23 35.805 ;
		RECT	2.18 35.215 2.23 35.345 ;
		RECT	2.18 32.795 2.23 32.925 ;
		RECT	2.18 32.335 2.23 32.465 ;
		RECT	2.18 29.915 2.23 30.045 ;
		RECT	2.18 29.455 2.23 29.585 ;
		RECT	2.18 27.035 2.23 27.165 ;
		RECT	2.18 26.575 2.23 26.705 ;
		RECT	2.18 24.155 2.23 24.285 ;
		RECT	2.18 23.695 2.23 23.825 ;
		RECT	2.18 21.275 2.23 21.405 ;
		RECT	2.18 20.815 2.23 20.945 ;
		RECT	2.18 18.395 2.23 18.525 ;
		RECT	2.18 17.935 2.23 18.065 ;
		RECT	2.18 15.515 2.23 15.645 ;
		RECT	2.18 15.055 2.23 15.185 ;
		RECT	2.18 12.635 2.23 12.765 ;
		RECT	2.18 170.575 2.23 170.705 ;
		RECT	2.18 168.155 2.23 168.285 ;
		RECT	2.18 12.175 2.23 12.305 ;
		RECT	2.18 9.755 2.23 9.885 ;
		RECT	2.18 9.295 2.23 9.425 ;
		RECT	2.18 6.875 2.23 7.005 ;
		RECT	2.18 6.415 2.23 6.545 ;
		RECT	2.18 3.995 2.23 4.125 ;
		RECT	2.18 3.535 2.23 3.665 ;
		RECT	2.18 1.115 2.23 1.245 ;
		RECT	2.18 167.695 2.23 167.825 ;
		RECT	2.18 165.275 2.23 165.405 ;
		RECT	2.18 164.815 2.23 164.945 ;
		RECT	2.18 162.395 2.23 162.525 ;
		RECT	2.18 161.935 2.23 162.065 ;
		RECT	2.18 159.515 2.23 159.645 ;
		RECT	2.18 159.055 2.23 159.185 ;
		RECT	2.18 156.635 2.23 156.765 ;
		RECT	1.38 184.975 1.43 185.105 ;
		RECT	4.51 184.975 4.56 185.105 ;
		RECT	3.06 184.515 3.11 184.645 ;
		RECT	1.405 182.555 1.455 182.685 ;
		RECT	4.51 182.555 4.56 182.685 ;
		RECT	1.38 156.175 1.43 156.305 ;
		RECT	4.51 156.175 4.56 156.305 ;
		RECT	3.06 155.715 3.11 155.845 ;
		RECT	1.405 153.755 1.455 153.885 ;
		RECT	4.51 153.755 4.56 153.885 ;
		RECT	1.38 153.295 1.43 153.425 ;
		RECT	4.51 153.295 4.56 153.425 ;
		RECT	3.06 152.835 3.11 152.965 ;
		RECT	1.405 150.875 1.455 151.005 ;
		RECT	4.51 150.875 4.56 151.005 ;
		RECT	1.38 150.415 1.43 150.545 ;
		RECT	4.51 150.415 4.56 150.545 ;
		RECT	3.06 149.955 3.11 150.085 ;
		RECT	1.405 147.995 1.455 148.125 ;
		RECT	4.51 147.995 4.56 148.125 ;
		RECT	1.38 147.535 1.43 147.665 ;
		RECT	4.51 147.535 4.56 147.665 ;
		RECT	3.06 147.075 3.11 147.205 ;
		RECT	1.405 145.115 1.455 145.245 ;
		RECT	4.51 145.115 4.56 145.245 ;
		RECT	1.38 144.655 1.43 144.785 ;
		RECT	4.51 144.655 4.56 144.785 ;
		RECT	3.06 144.195 3.11 144.325 ;
		RECT	1.405 142.235 1.455 142.365 ;
		RECT	4.51 142.235 4.56 142.365 ;
		RECT	1.38 141.775 1.43 141.905 ;
		RECT	4.51 141.775 4.56 141.905 ;
		RECT	3.06 141.315 3.11 141.445 ;
		RECT	1.405 139.355 1.455 139.485 ;
		RECT	4.51 139.355 4.56 139.485 ;
		RECT	1.38 138.895 1.43 139.025 ;
		RECT	4.51 138.895 4.56 139.025 ;
		RECT	3.06 138.435 3.11 138.565 ;
		RECT	1.405 136.475 1.455 136.605 ;
		RECT	4.51 136.475 4.56 136.605 ;
		RECT	1.38 136.015 1.43 136.145 ;
		RECT	4.51 136.015 4.56 136.145 ;
		RECT	3.06 135.555 3.11 135.685 ;
		RECT	1.405 133.595 1.455 133.725 ;
		RECT	4.51 133.595 4.56 133.725 ;
		RECT	1.38 133.135 1.43 133.265 ;
		RECT	4.51 133.135 4.56 133.265 ;
		RECT	3.06 132.675 3.11 132.805 ;
		RECT	1.405 130.715 1.455 130.845 ;
		RECT	4.51 130.715 4.56 130.845 ;
		RECT	1.38 130.255 1.43 130.385 ;
		RECT	4.51 130.255 4.56 130.385 ;
		RECT	3.06 129.795 3.11 129.925 ;
		RECT	1.405 127.835 1.455 127.965 ;
		RECT	4.51 127.835 4.56 127.965 ;
		RECT	1.38 182.095 1.43 182.225 ;
		RECT	4.51 182.095 4.56 182.225 ;
		RECT	3.06 181.635 3.11 181.765 ;
		RECT	1.405 179.675 1.455 179.805 ;
		RECT	4.51 179.675 4.56 179.805 ;
		RECT	1.38 127.375 1.43 127.505 ;
		RECT	4.51 127.375 4.56 127.505 ;
		RECT	3.06 126.915 3.11 127.045 ;
		RECT	1.405 124.955 1.455 125.085 ;
		RECT	4.51 124.955 4.56 125.085 ;
		RECT	1.38 124.495 1.43 124.625 ;
		RECT	4.51 124.495 4.56 124.625 ;
		RECT	3.06 124.035 3.11 124.165 ;
		RECT	1.405 122.075 1.455 122.205 ;
		RECT	4.51 122.075 4.56 122.205 ;
		RECT	1.38 121.615 1.43 121.745 ;
		RECT	4.51 121.615 4.56 121.745 ;
		RECT	3.06 121.155 3.11 121.285 ;
		RECT	1.405 119.195 1.455 119.325 ;
		RECT	4.51 119.195 4.56 119.325 ;
		RECT	1.38 118.735 1.43 118.865 ;
		RECT	4.51 118.735 4.56 118.865 ;
		RECT	3.06 118.275 3.11 118.405 ;
		RECT	1.405 116.315 1.455 116.445 ;
		RECT	4.51 116.315 4.56 116.445 ;
		RECT	1.38 115.855 1.43 115.985 ;
		RECT	4.51 115.855 4.56 115.985 ;
		RECT	3.06 115.395 3.11 115.525 ;
		RECT	1.405 113.435 1.455 113.565 ;
		RECT	4.51 113.435 4.56 113.565 ;
		RECT	1.38 112.975 1.43 113.105 ;
		RECT	4.51 112.975 4.56 113.105 ;
		RECT	3.06 112.515 3.11 112.645 ;
		RECT	1.405 110.555 1.455 110.685 ;
		RECT	4.51 110.555 4.56 110.685 ;
		RECT	1.38 110.095 1.43 110.225 ;
		RECT	4.51 110.095 4.56 110.225 ;
		RECT	3.06 109.635 3.11 109.765 ;
		RECT	1.405 107.675 1.455 107.805 ;
		RECT	4.51 107.675 4.56 107.805 ;
		RECT	1.38 107.215 1.43 107.345 ;
		RECT	4.51 107.215 4.56 107.345 ;
		RECT	3.06 106.755 3.11 106.885 ;
		RECT	1.405 104.795 1.455 104.925 ;
		RECT	4.51 104.795 4.56 104.925 ;
		RECT	1.38 104.335 1.43 104.465 ;
		RECT	4.51 104.335 4.56 104.465 ;
		RECT	3.06 103.875 3.11 104.005 ;
		RECT	1.405 101.915 1.455 102.045 ;
		RECT	4.51 101.915 4.56 102.045 ;
		RECT	1.38 101.455 1.43 101.585 ;
		RECT	4.51 101.455 4.56 101.585 ;
		RECT	3.06 100.995 3.11 101.125 ;
		RECT	1.405 99.035 1.455 99.165 ;
		RECT	4.51 99.035 4.56 99.165 ;
		RECT	1.38 179.215 1.43 179.345 ;
		RECT	4.51 179.215 4.56 179.345 ;
		RECT	3.06 178.755 3.11 178.885 ;
		RECT	1.405 176.795 1.455 176.925 ;
		RECT	4.51 176.795 4.56 176.925 ;
		RECT	1.38 98.575 1.43 98.705 ;
		RECT	4.51 98.575 4.56 98.705 ;
		RECT	3.06 98.115 3.11 98.245 ;
		RECT	1.405 96.155 1.455 96.285 ;
		RECT	4.51 96.155 4.56 96.285 ;
		RECT	1.38 95.695 1.43 95.825 ;
		RECT	4.51 95.695 4.56 95.825 ;
		RECT	3.06 95.235 3.11 95.365 ;
		RECT	1.405 93.275 1.455 93.405 ;
		RECT	4.51 93.275 4.56 93.405 ;
		RECT	1.38 92.815 1.43 92.945 ;
		RECT	4.51 92.815 4.56 92.945 ;
		RECT	3.06 92.355 3.11 92.485 ;
		RECT	1.405 90.395 1.455 90.525 ;
		RECT	4.51 90.395 4.56 90.525 ;
		RECT	1.38 89.935 1.43 90.065 ;
		RECT	4.51 89.935 4.56 90.065 ;
		RECT	3.06 89.475 3.11 89.605 ;
		RECT	1.405 87.515 1.455 87.645 ;
		RECT	4.51 87.515 4.56 87.645 ;
		RECT	1.38 87.055 1.43 87.185 ;
		RECT	4.51 87.055 4.56 87.185 ;
		RECT	3.06 86.595 3.11 86.725 ;
		RECT	1.405 84.635 1.455 84.765 ;
		RECT	4.51 84.635 4.56 84.765 ;
		RECT	1.38 84.175 1.43 84.305 ;
		RECT	4.51 84.175 4.56 84.305 ;
		RECT	3.06 83.715 3.11 83.845 ;
		RECT	1.405 81.755 1.455 81.885 ;
		RECT	4.51 81.755 4.56 81.885 ;
		RECT	1.38 81.295 1.43 81.425 ;
		RECT	4.51 81.295 4.56 81.425 ;
		RECT	3.06 80.835 3.11 80.965 ;
		RECT	1.405 78.875 1.455 79.005 ;
		RECT	4.51 78.875 4.56 79.005 ;
		RECT	1.38 78.415 1.43 78.545 ;
		RECT	4.51 78.415 4.56 78.545 ;
		RECT	3.06 77.955 3.11 78.085 ;
		RECT	1.405 75.995 1.455 76.125 ;
		RECT	4.51 75.995 4.56 76.125 ;
		RECT	1.38 75.535 1.43 75.665 ;
		RECT	4.51 75.535 4.56 75.665 ;
		RECT	3.06 75.075 3.11 75.205 ;
		RECT	1.405 73.115 1.455 73.245 ;
		RECT	4.51 73.115 4.56 73.245 ;
		RECT	1.38 72.655 1.43 72.785 ;
		RECT	4.51 72.655 4.56 72.785 ;
		RECT	3.06 72.195 3.11 72.325 ;
		RECT	1.405 70.235 1.455 70.365 ;
		RECT	4.51 70.235 4.56 70.365 ;
		RECT	1.38 176.335 1.43 176.465 ;
		RECT	4.51 176.335 4.56 176.465 ;
		RECT	3.06 175.875 3.11 176.005 ;
		RECT	1.405 173.915 1.455 174.045 ;
		RECT	4.51 173.915 4.56 174.045 ;
		RECT	1.38 69.775 1.43 69.905 ;
		RECT	4.51 69.775 4.56 69.905 ;
		RECT	3.06 69.315 3.11 69.445 ;
		RECT	1.405 67.355 1.455 67.485 ;
		RECT	4.51 67.355 4.56 67.485 ;
		RECT	1.38 66.895 1.43 67.025 ;
		RECT	4.51 66.895 4.56 67.025 ;
		RECT	3.06 66.435 3.11 66.565 ;
		RECT	1.405 64.475 1.455 64.605 ;
		RECT	4.51 64.475 4.56 64.605 ;
		RECT	1.38 64.015 1.43 64.145 ;
		RECT	4.51 64.015 4.56 64.145 ;
		RECT	3.06 63.555 3.11 63.685 ;
		RECT	1.405 61.595 1.455 61.725 ;
		RECT	4.51 61.595 4.56 61.725 ;
		RECT	1.38 61.135 1.43 61.265 ;
		RECT	4.51 61.135 4.56 61.265 ;
		RECT	3.06 60.675 3.11 60.805 ;
		RECT	1.405 58.715 1.455 58.845 ;
		RECT	4.51 58.715 4.56 58.845 ;
		RECT	1.38 58.255 1.43 58.385 ;
		RECT	4.51 58.255 4.56 58.385 ;
		RECT	3.06 57.795 3.11 57.925 ;
		RECT	1.405 55.835 1.455 55.965 ;
		RECT	4.51 55.835 4.56 55.965 ;
		RECT	1.38 55.375 1.43 55.505 ;
		RECT	4.51 55.375 4.56 55.505 ;
		RECT	3.06 54.915 3.11 55.045 ;
		RECT	1.405 52.955 1.455 53.085 ;
		RECT	4.51 52.955 4.56 53.085 ;
		RECT	1.38 52.495 1.43 52.625 ;
		RECT	4.51 52.495 4.56 52.625 ;
		RECT	3.06 52.035 3.11 52.165 ;
		RECT	1.405 50.075 1.455 50.205 ;
		RECT	4.51 50.075 4.56 50.205 ;
		RECT	1.38 49.615 1.43 49.745 ;
		RECT	4.51 49.615 4.56 49.745 ;
		RECT	3.06 49.155 3.11 49.285 ;
		RECT	1.405 47.195 1.455 47.325 ;
		RECT	4.51 47.195 4.56 47.325 ;
		RECT	1.38 46.735 1.43 46.865 ;
		RECT	4.51 46.735 4.56 46.865 ;
		RECT	3.06 46.275 3.11 46.405 ;
		RECT	1.405 44.315 1.455 44.445 ;
		RECT	4.51 44.315 4.56 44.445 ;
		RECT	1.38 43.855 1.43 43.985 ;
		RECT	4.51 43.855 4.56 43.985 ;
		RECT	3.06 43.395 3.11 43.525 ;
		RECT	1.405 41.435 1.455 41.565 ;
		RECT	4.51 41.435 4.56 41.565 ;
		RECT	1.38 173.455 1.43 173.585 ;
		RECT	4.51 173.455 4.56 173.585 ;
		RECT	3.06 172.995 3.11 173.125 ;
		RECT	1.405 171.035 1.455 171.165 ;
		RECT	4.51 171.035 4.56 171.165 ;
		RECT	1.38 40.975 1.43 41.105 ;
		RECT	4.51 40.975 4.56 41.105 ;
		RECT	3.06 40.515 3.11 40.645 ;
		RECT	1.405 38.555 1.455 38.685 ;
		RECT	4.51 38.555 4.56 38.685 ;
		RECT	1.38 38.095 1.43 38.225 ;
		RECT	4.51 38.095 4.56 38.225 ;
		RECT	3.06 37.635 3.11 37.765 ;
		RECT	1.405 35.675 1.455 35.805 ;
		RECT	4.51 35.675 4.56 35.805 ;
		RECT	1.38 35.215 1.43 35.345 ;
		RECT	4.51 35.215 4.56 35.345 ;
		RECT	3.06 34.755 3.11 34.885 ;
		RECT	1.405 32.795 1.455 32.925 ;
		RECT	4.51 32.795 4.56 32.925 ;
		RECT	1.38 32.335 1.43 32.465 ;
		RECT	4.51 32.335 4.56 32.465 ;
		RECT	3.06 31.875 3.11 32.005 ;
		RECT	1.405 29.915 1.455 30.045 ;
		RECT	4.51 29.915 4.56 30.045 ;
		RECT	1.38 29.455 1.43 29.585 ;
		RECT	4.51 29.455 4.56 29.585 ;
		RECT	3.06 28.995 3.11 29.125 ;
		RECT	1.405 27.035 1.455 27.165 ;
		RECT	4.51 27.035 4.56 27.165 ;
		RECT	1.38 26.575 1.43 26.705 ;
		RECT	4.51 26.575 4.56 26.705 ;
		RECT	3.06 26.115 3.11 26.245 ;
		RECT	1.405 24.155 1.455 24.285 ;
		RECT	4.51 24.155 4.56 24.285 ;
		RECT	1.38 23.695 1.43 23.825 ;
		RECT	4.51 23.695 4.56 23.825 ;
		RECT	3.06 23.235 3.11 23.365 ;
		RECT	1.405 21.275 1.455 21.405 ;
		RECT	4.51 21.275 4.56 21.405 ;
		RECT	1.38 20.815 1.43 20.945 ;
		RECT	4.51 20.815 4.56 20.945 ;
		RECT	3.06 20.355 3.11 20.485 ;
		RECT	1.405 18.395 1.455 18.525 ;
		RECT	4.51 18.395 4.56 18.525 ;
		RECT	1.38 17.935 1.43 18.065 ;
		RECT	4.51 17.935 4.56 18.065 ;
		RECT	3.06 17.475 3.11 17.605 ;
		RECT	1.405 15.515 1.455 15.645 ;
		RECT	4.51 15.515 4.56 15.645 ;
		RECT	1.38 15.055 1.43 15.185 ;
		RECT	4.51 15.055 4.56 15.185 ;
		RECT	3.06 14.595 3.11 14.725 ;
		RECT	1.405 12.635 1.455 12.765 ;
		RECT	4.51 12.635 4.56 12.765 ;
		RECT	1.38 170.575 1.43 170.705 ;
		RECT	4.51 170.575 4.56 170.705 ;
		RECT	3.06 170.115 3.11 170.245 ;
		RECT	1.405 168.155 1.455 168.285 ;
		RECT	4.51 168.155 4.56 168.285 ;
		RECT	1.38 12.175 1.43 12.305 ;
		RECT	4.51 12.175 4.56 12.305 ;
		RECT	3.06 11.715 3.11 11.845 ;
		RECT	1.405 9.755 1.455 9.885 ;
		RECT	4.51 9.755 4.56 9.885 ;
		RECT	1.38 9.295 1.43 9.425 ;
		RECT	4.51 9.295 4.56 9.425 ;
		RECT	3.06 8.835 3.11 8.965 ;
		RECT	1.405 6.875 1.455 7.005 ;
		RECT	4.51 6.875 4.56 7.005 ;
		RECT	1.38 6.415 1.43 6.545 ;
		RECT	4.51 6.415 4.56 6.545 ;
		RECT	3.06 5.955 3.11 6.085 ;
		RECT	1.405 3.995 1.455 4.125 ;
		RECT	4.51 3.995 4.56 4.125 ;
		RECT	1.38 3.535 1.43 3.665 ;
		RECT	4.51 3.535 4.56 3.665 ;
		RECT	3.06 3.075 3.11 3.205 ;
		RECT	1.405 1.115 1.455 1.245 ;
		RECT	4.51 1.115 4.56 1.245 ;
		RECT	1.38 167.695 1.43 167.825 ;
		RECT	4.51 167.695 4.56 167.825 ;
		RECT	3.06 167.235 3.11 167.365 ;
		RECT	1.405 165.275 1.455 165.405 ;
		RECT	4.51 165.275 4.56 165.405 ;
		RECT	1.38 164.815 1.43 164.945 ;
		RECT	4.51 164.815 4.56 164.945 ;
		RECT	3.06 164.355 3.11 164.485 ;
		RECT	1.405 162.395 1.455 162.525 ;
		RECT	4.51 162.395 4.56 162.525 ;
		RECT	1.38 161.935 1.43 162.065 ;
		RECT	4.51 161.935 4.56 162.065 ;
		RECT	3.06 161.475 3.11 161.605 ;
		RECT	1.405 159.515 1.455 159.645 ;
		RECT	4.51 159.515 4.56 159.645 ;
		RECT	1.38 159.055 1.43 159.185 ;
		RECT	4.51 159.055 4.56 159.185 ;
		RECT	3.06 158.595 3.11 158.725 ;
		RECT	1.405 156.635 1.455 156.765 ;
		RECT	4.51 156.635 4.56 156.765 ;
		RECT	3.06 182.095 3.11 182.225 ;
		RECT	1.085 181.635 1.135 181.765 ;
		RECT	1.405 181.675 1.455 181.725 ;
		RECT	4.47 181.675 4.6 181.725 ;
		RECT	3.06 179.675 3.11 179.805 ;
		RECT	1.57 179.445 1.62 179.575 ;
		RECT	2.58 179.445 2.63 179.575 ;
		RECT	3.84 179.445 3.89 179.575 ;
		RECT	5.675 179.445 5.725 179.575 ;
		RECT	3.06 156.175 3.11 156.305 ;
		RECT	1.085 155.715 1.135 155.845 ;
		RECT	1.405 155.755 1.455 155.805 ;
		RECT	4.47 155.755 4.6 155.805 ;
		RECT	3.06 153.755 3.11 153.885 ;
		RECT	1.57 153.525 1.62 153.655 ;
		RECT	2.58 153.525 2.63 153.655 ;
		RECT	3.84 153.525 3.89 153.655 ;
		RECT	5.675 153.525 5.725 153.655 ;
		RECT	3.06 153.295 3.11 153.425 ;
		RECT	1.085 152.835 1.135 152.965 ;
		RECT	1.405 152.875 1.455 152.925 ;
		RECT	4.47 152.875 4.6 152.925 ;
		RECT	3.06 150.875 3.11 151.005 ;
		RECT	1.57 150.645 1.62 150.775 ;
		RECT	2.58 150.645 2.63 150.775 ;
		RECT	3.84 150.645 3.89 150.775 ;
		RECT	5.675 150.645 5.725 150.775 ;
		RECT	3.06 150.415 3.11 150.545 ;
		RECT	1.085 149.955 1.135 150.085 ;
		RECT	1.405 149.995 1.455 150.045 ;
		RECT	4.47 149.995 4.6 150.045 ;
		RECT	3.06 147.995 3.11 148.125 ;
		RECT	1.57 147.765 1.62 147.895 ;
		RECT	2.58 147.765 2.63 147.895 ;
		RECT	3.84 147.765 3.89 147.895 ;
		RECT	5.675 147.765 5.725 147.895 ;
		RECT	3.06 147.535 3.11 147.665 ;
		RECT	1.085 147.075 1.135 147.205 ;
		RECT	1.405 147.115 1.455 147.165 ;
		RECT	4.47 147.115 4.6 147.165 ;
		RECT	3.06 145.115 3.11 145.245 ;
		RECT	1.57 144.885 1.62 145.015 ;
		RECT	2.58 144.885 2.63 145.015 ;
		RECT	3.84 144.885 3.89 145.015 ;
		RECT	5.675 144.885 5.725 145.015 ;
		RECT	3.06 144.655 3.11 144.785 ;
		RECT	1.085 144.195 1.135 144.325 ;
		RECT	1.405 144.235 1.455 144.285 ;
		RECT	4.47 144.235 4.6 144.285 ;
		RECT	3.06 142.235 3.11 142.365 ;
		RECT	1.57 142.005 1.62 142.135 ;
		RECT	2.58 142.005 2.63 142.135 ;
		RECT	3.84 142.005 3.89 142.135 ;
		RECT	5.675 142.005 5.725 142.135 ;
		RECT	3.06 141.775 3.11 141.905 ;
		RECT	1.085 141.315 1.135 141.445 ;
		RECT	1.405 141.355 1.455 141.405 ;
		RECT	4.47 141.355 4.6 141.405 ;
		RECT	3.06 139.355 3.11 139.485 ;
		RECT	1.57 139.125 1.62 139.255 ;
		RECT	2.58 139.125 2.63 139.255 ;
		RECT	3.84 139.125 3.89 139.255 ;
		RECT	5.675 139.125 5.725 139.255 ;
		RECT	3.06 138.895 3.11 139.025 ;
		RECT	1.085 138.435 1.135 138.565 ;
		RECT	1.405 138.475 1.455 138.525 ;
		RECT	4.47 138.475 4.6 138.525 ;
		RECT	3.06 136.475 3.11 136.605 ;
		RECT	1.57 136.245 1.62 136.375 ;
		RECT	2.58 136.245 2.63 136.375 ;
		RECT	3.84 136.245 3.89 136.375 ;
		RECT	5.675 136.245 5.725 136.375 ;
		RECT	3.06 136.015 3.11 136.145 ;
		RECT	1.085 135.555 1.135 135.685 ;
		RECT	1.405 135.595 1.455 135.645 ;
		RECT	4.47 135.595 4.6 135.645 ;
		RECT	3.06 133.595 3.11 133.725 ;
		RECT	1.57 133.365 1.62 133.495 ;
		RECT	2.58 133.365 2.63 133.495 ;
		RECT	3.84 133.365 3.89 133.495 ;
		RECT	5.675 133.365 5.725 133.495 ;
		RECT	3.06 133.135 3.11 133.265 ;
		RECT	1.085 132.675 1.135 132.805 ;
		RECT	1.405 132.715 1.455 132.765 ;
		RECT	4.47 132.715 4.6 132.765 ;
		RECT	3.06 130.715 3.11 130.845 ;
		RECT	1.57 130.485 1.62 130.615 ;
		RECT	2.58 130.485 2.63 130.615 ;
		RECT	3.84 130.485 3.89 130.615 ;
		RECT	5.675 130.485 5.725 130.615 ;
		RECT	3.06 130.255 3.11 130.385 ;
		RECT	1.085 129.795 1.135 129.925 ;
		RECT	1.405 129.835 1.455 129.885 ;
		RECT	4.47 129.835 4.6 129.885 ;
		RECT	3.06 127.835 3.11 127.965 ;
		RECT	1.57 127.605 1.62 127.735 ;
		RECT	2.58 127.605 2.63 127.735 ;
		RECT	3.84 127.605 3.89 127.735 ;
		RECT	5.675 127.605 5.725 127.735 ;
		RECT	3.06 179.215 3.11 179.345 ;
		RECT	1.085 178.755 1.135 178.885 ;
		RECT	1.405 178.795 1.455 178.845 ;
		RECT	4.47 178.795 4.6 178.845 ;
		RECT	3.06 176.795 3.11 176.925 ;
		RECT	1.57 176.565 1.62 176.695 ;
		RECT	2.58 176.565 2.63 176.695 ;
		RECT	3.84 176.565 3.89 176.695 ;
		RECT	5.675 176.565 5.725 176.695 ;
		RECT	3.06 127.375 3.11 127.505 ;
		RECT	1.085 126.915 1.135 127.045 ;
		RECT	1.405 126.955 1.455 127.005 ;
		RECT	4.47 126.955 4.6 127.005 ;
		RECT	3.06 124.955 3.11 125.085 ;
		RECT	1.57 124.725 1.62 124.855 ;
		RECT	2.58 124.725 2.63 124.855 ;
		RECT	3.84 124.725 3.89 124.855 ;
		RECT	5.675 124.725 5.725 124.855 ;
		RECT	3.06 124.495 3.11 124.625 ;
		RECT	1.085 124.035 1.135 124.165 ;
		RECT	1.405 124.075 1.455 124.125 ;
		RECT	4.47 124.075 4.6 124.125 ;
		RECT	3.06 122.075 3.11 122.205 ;
		RECT	1.57 121.845 1.62 121.975 ;
		RECT	2.58 121.845 2.63 121.975 ;
		RECT	3.84 121.845 3.89 121.975 ;
		RECT	5.675 121.845 5.725 121.975 ;
		RECT	3.06 121.615 3.11 121.745 ;
		RECT	1.085 121.155 1.135 121.285 ;
		RECT	1.405 121.195 1.455 121.245 ;
		RECT	4.47 121.195 4.6 121.245 ;
		RECT	3.06 119.195 3.11 119.325 ;
		RECT	1.57 118.965 1.62 119.095 ;
		RECT	2.58 118.965 2.63 119.095 ;
		RECT	3.84 118.965 3.89 119.095 ;
		RECT	5.675 118.965 5.725 119.095 ;
		RECT	3.06 118.735 3.11 118.865 ;
		RECT	1.085 118.275 1.135 118.405 ;
		RECT	1.405 118.315 1.455 118.365 ;
		RECT	4.47 118.315 4.6 118.365 ;
		RECT	3.06 116.315 3.11 116.445 ;
		RECT	1.57 116.085 1.62 116.215 ;
		RECT	2.58 116.085 2.63 116.215 ;
		RECT	3.84 116.085 3.89 116.215 ;
		RECT	5.675 116.085 5.725 116.215 ;
		RECT	3.06 115.855 3.11 115.985 ;
		RECT	1.085 115.395 1.135 115.525 ;
		RECT	1.405 115.435 1.455 115.485 ;
		RECT	4.47 115.435 4.6 115.485 ;
		RECT	3.06 113.435 3.11 113.565 ;
		RECT	1.57 113.205 1.62 113.335 ;
		RECT	2.58 113.205 2.63 113.335 ;
		RECT	3.84 113.205 3.89 113.335 ;
		RECT	5.675 113.205 5.725 113.335 ;
		RECT	3.06 112.975 3.11 113.105 ;
		RECT	1.085 112.515 1.135 112.645 ;
		RECT	1.405 112.555 1.455 112.605 ;
		RECT	4.47 112.555 4.6 112.605 ;
		RECT	3.06 110.555 3.11 110.685 ;
		RECT	1.57 110.325 1.62 110.455 ;
		RECT	2.58 110.325 2.63 110.455 ;
		RECT	3.84 110.325 3.89 110.455 ;
		RECT	5.675 110.325 5.725 110.455 ;
		RECT	3.06 110.095 3.11 110.225 ;
		RECT	1.085 109.635 1.135 109.765 ;
		RECT	1.405 109.675 1.455 109.725 ;
		RECT	4.47 109.675 4.6 109.725 ;
		RECT	3.06 107.675 3.11 107.805 ;
		RECT	1.57 107.445 1.62 107.575 ;
		RECT	2.58 107.445 2.63 107.575 ;
		RECT	3.84 107.445 3.89 107.575 ;
		RECT	5.675 107.445 5.725 107.575 ;
		RECT	3.06 107.215 3.11 107.345 ;
		RECT	1.085 106.755 1.135 106.885 ;
		RECT	1.405 106.795 1.455 106.845 ;
		RECT	4.47 106.795 4.6 106.845 ;
		RECT	3.06 104.795 3.11 104.925 ;
		RECT	1.57 104.565 1.62 104.695 ;
		RECT	2.58 104.565 2.63 104.695 ;
		RECT	3.84 104.565 3.89 104.695 ;
		RECT	5.675 104.565 5.725 104.695 ;
		RECT	3.06 104.335 3.11 104.465 ;
		RECT	1.085 103.875 1.135 104.005 ;
		RECT	1.405 103.915 1.455 103.965 ;
		RECT	4.47 103.915 4.6 103.965 ;
		RECT	3.06 101.915 3.11 102.045 ;
		RECT	1.57 101.685 1.62 101.815 ;
		RECT	2.58 101.685 2.63 101.815 ;
		RECT	3.84 101.685 3.89 101.815 ;
		RECT	5.675 101.685 5.725 101.815 ;
		RECT	3.06 101.455 3.11 101.585 ;
		RECT	1.085 100.995 1.135 101.125 ;
		RECT	1.405 101.035 1.455 101.085 ;
		RECT	4.47 101.035 4.6 101.085 ;
		RECT	3.06 99.035 3.11 99.165 ;
		RECT	1.57 98.805 1.62 98.935 ;
		RECT	2.58 98.805 2.63 98.935 ;
		RECT	3.84 98.805 3.89 98.935 ;
		RECT	5.675 98.805 5.725 98.935 ;
		RECT	3.06 176.335 3.11 176.465 ;
		RECT	1.085 175.875 1.135 176.005 ;
		RECT	1.405 175.915 1.455 175.965 ;
		RECT	4.47 175.915 4.6 175.965 ;
		RECT	3.06 173.915 3.11 174.045 ;
		RECT	1.57 173.685 1.62 173.815 ;
		RECT	2.58 173.685 2.63 173.815 ;
		RECT	3.84 173.685 3.89 173.815 ;
		RECT	5.675 173.685 5.725 173.815 ;
		RECT	3.06 98.575 3.11 98.705 ;
		RECT	1.085 98.115 1.135 98.245 ;
		RECT	1.405 98.155 1.455 98.205 ;
		RECT	4.47 98.155 4.6 98.205 ;
		RECT	3.06 96.155 3.11 96.285 ;
		RECT	1.57 95.925 1.62 96.055 ;
		RECT	2.58 95.925 2.63 96.055 ;
		RECT	3.84 95.925 3.89 96.055 ;
		RECT	5.675 95.925 5.725 96.055 ;
		RECT	3.06 95.695 3.11 95.825 ;
		RECT	1.085 95.235 1.135 95.365 ;
		RECT	1.405 95.275 1.455 95.325 ;
		RECT	4.47 95.275 4.6 95.325 ;
		RECT	3.06 93.275 3.11 93.405 ;
		RECT	1.57 93.045 1.62 93.175 ;
		RECT	2.58 93.045 2.63 93.175 ;
		RECT	3.84 93.045 3.89 93.175 ;
		RECT	5.675 93.045 5.725 93.175 ;
		RECT	3.06 92.815 3.11 92.945 ;
		RECT	1.085 92.355 1.135 92.485 ;
		RECT	1.405 92.395 1.455 92.445 ;
		RECT	4.47 92.395 4.6 92.445 ;
		RECT	3.06 90.395 3.11 90.525 ;
		RECT	1.57 90.165 1.62 90.295 ;
		RECT	2.58 90.165 2.63 90.295 ;
		RECT	3.84 90.165 3.89 90.295 ;
		RECT	5.675 90.165 5.725 90.295 ;
		RECT	3.06 89.935 3.11 90.065 ;
		RECT	1.085 89.475 1.135 89.605 ;
		RECT	1.405 89.515 1.455 89.565 ;
		RECT	4.47 89.515 4.6 89.565 ;
		RECT	3.06 87.515 3.11 87.645 ;
		RECT	1.57 87.285 1.62 87.415 ;
		RECT	2.58 87.285 2.63 87.415 ;
		RECT	3.84 87.285 3.89 87.415 ;
		RECT	5.675 87.285 5.725 87.415 ;
		RECT	3.06 87.055 3.11 87.185 ;
		RECT	1.085 86.595 1.135 86.725 ;
		RECT	1.405 86.635 1.455 86.685 ;
		RECT	4.47 86.635 4.6 86.685 ;
		RECT	3.06 84.635 3.11 84.765 ;
		RECT	1.57 84.405 1.62 84.535 ;
		RECT	2.58 84.405 2.63 84.535 ;
		RECT	3.84 84.405 3.89 84.535 ;
		RECT	5.675 84.405 5.725 84.535 ;
		RECT	3.06 84.175 3.11 84.305 ;
		RECT	1.085 83.715 1.135 83.845 ;
		RECT	1.405 83.755 1.455 83.805 ;
		RECT	4.47 83.755 4.6 83.805 ;
		RECT	3.06 81.755 3.11 81.885 ;
		RECT	1.57 81.525 1.62 81.655 ;
		RECT	2.58 81.525 2.63 81.655 ;
		RECT	3.84 81.525 3.89 81.655 ;
		RECT	5.675 81.525 5.725 81.655 ;
		RECT	3.06 81.295 3.11 81.425 ;
		RECT	1.085 80.835 1.135 80.965 ;
		RECT	1.405 80.875 1.455 80.925 ;
		RECT	4.47 80.875 4.6 80.925 ;
		RECT	3.06 78.875 3.11 79.005 ;
		RECT	1.57 78.645 1.62 78.775 ;
		RECT	2.58 78.645 2.63 78.775 ;
		RECT	3.84 78.645 3.89 78.775 ;
		RECT	5.675 78.645 5.725 78.775 ;
		RECT	3.06 78.415 3.11 78.545 ;
		RECT	1.085 77.955 1.135 78.085 ;
		RECT	1.405 77.995 1.455 78.045 ;
		RECT	4.47 77.995 4.6 78.045 ;
		RECT	3.06 75.995 3.11 76.125 ;
		RECT	1.57 75.765 1.62 75.895 ;
		RECT	2.58 75.765 2.63 75.895 ;
		RECT	3.84 75.765 3.89 75.895 ;
		RECT	5.675 75.765 5.725 75.895 ;
		RECT	3.06 75.535 3.11 75.665 ;
		RECT	1.085 75.075 1.135 75.205 ;
		RECT	1.405 75.115 1.455 75.165 ;
		RECT	4.47 75.115 4.6 75.165 ;
		RECT	3.06 73.115 3.11 73.245 ;
		RECT	1.57 72.885 1.62 73.015 ;
		RECT	2.58 72.885 2.63 73.015 ;
		RECT	3.84 72.885 3.89 73.015 ;
		RECT	5.675 72.885 5.725 73.015 ;
		RECT	3.06 72.655 3.11 72.785 ;
		RECT	1.085 72.195 1.135 72.325 ;
		RECT	1.405 72.235 1.455 72.285 ;
		RECT	4.47 72.235 4.6 72.285 ;
		RECT	3.06 70.235 3.11 70.365 ;
		RECT	1.57 70.005 1.62 70.135 ;
		RECT	2.58 70.005 2.63 70.135 ;
		RECT	3.84 70.005 3.89 70.135 ;
		RECT	5.675 70.005 5.725 70.135 ;
		RECT	3.06 173.455 3.11 173.585 ;
		RECT	1.085 172.995 1.135 173.125 ;
		RECT	1.405 173.035 1.455 173.085 ;
		RECT	4.47 173.035 4.6 173.085 ;
		RECT	3.06 171.035 3.11 171.165 ;
		RECT	1.57 170.805 1.62 170.935 ;
		RECT	2.58 170.805 2.63 170.935 ;
		RECT	3.84 170.805 3.89 170.935 ;
		RECT	5.675 170.805 5.725 170.935 ;
		RECT	3.06 69.775 3.11 69.905 ;
		RECT	1.085 69.315 1.135 69.445 ;
		RECT	1.405 69.355 1.455 69.405 ;
		RECT	4.47 69.355 4.6 69.405 ;
		RECT	3.06 67.355 3.11 67.485 ;
		RECT	1.57 67.125 1.62 67.255 ;
		RECT	2.58 67.125 2.63 67.255 ;
		RECT	3.84 67.125 3.89 67.255 ;
		RECT	5.675 67.125 5.725 67.255 ;
		RECT	3.06 66.895 3.11 67.025 ;
		RECT	1.085 66.435 1.135 66.565 ;
		RECT	1.405 66.475 1.455 66.525 ;
		RECT	4.47 66.475 4.6 66.525 ;
		RECT	3.06 64.475 3.11 64.605 ;
		RECT	1.57 64.245 1.62 64.375 ;
		RECT	2.58 64.245 2.63 64.375 ;
		RECT	3.84 64.245 3.89 64.375 ;
		RECT	5.675 64.245 5.725 64.375 ;
		RECT	3.06 64.015 3.11 64.145 ;
		RECT	1.085 63.555 1.135 63.685 ;
		RECT	1.405 63.595 1.455 63.645 ;
		RECT	4.47 63.595 4.6 63.645 ;
		RECT	3.06 61.595 3.11 61.725 ;
		RECT	1.57 61.365 1.62 61.495 ;
		RECT	2.58 61.365 2.63 61.495 ;
		RECT	3.84 61.365 3.89 61.495 ;
		RECT	5.675 61.365 5.725 61.495 ;
		RECT	3.06 61.135 3.11 61.265 ;
		RECT	1.085 60.675 1.135 60.805 ;
		RECT	1.405 60.715 1.455 60.765 ;
		RECT	4.47 60.715 4.6 60.765 ;
		RECT	3.06 58.715 3.11 58.845 ;
		RECT	1.57 58.485 1.62 58.615 ;
		RECT	2.58 58.485 2.63 58.615 ;
		RECT	3.84 58.485 3.89 58.615 ;
		RECT	5.675 58.485 5.725 58.615 ;
		RECT	3.06 58.255 3.11 58.385 ;
		RECT	1.085 57.795 1.135 57.925 ;
		RECT	1.405 57.835 1.455 57.885 ;
		RECT	4.47 57.835 4.6 57.885 ;
		RECT	3.06 55.835 3.11 55.965 ;
		RECT	1.57 55.605 1.62 55.735 ;
		RECT	2.58 55.605 2.63 55.735 ;
		RECT	3.84 55.605 3.89 55.735 ;
		RECT	5.675 55.605 5.725 55.735 ;
		RECT	3.06 55.375 3.11 55.505 ;
		RECT	1.085 54.915 1.135 55.045 ;
		RECT	1.405 54.955 1.455 55.005 ;
		RECT	4.47 54.955 4.6 55.005 ;
		RECT	3.06 52.955 3.11 53.085 ;
		RECT	1.57 52.725 1.62 52.855 ;
		RECT	2.58 52.725 2.63 52.855 ;
		RECT	3.84 52.725 3.89 52.855 ;
		RECT	5.675 52.725 5.725 52.855 ;
		RECT	3.06 52.495 3.11 52.625 ;
		RECT	1.085 52.035 1.135 52.165 ;
		RECT	1.405 52.075 1.455 52.125 ;
		RECT	4.47 52.075 4.6 52.125 ;
		RECT	3.06 50.075 3.11 50.205 ;
		RECT	1.57 49.845 1.62 49.975 ;
		RECT	2.58 49.845 2.63 49.975 ;
		RECT	3.84 49.845 3.89 49.975 ;
		RECT	5.675 49.845 5.725 49.975 ;
		RECT	3.06 49.615 3.11 49.745 ;
		RECT	1.085 49.155 1.135 49.285 ;
		RECT	1.405 49.195 1.455 49.245 ;
		RECT	4.47 49.195 4.6 49.245 ;
		RECT	3.06 47.195 3.11 47.325 ;
		RECT	1.57 46.965 1.62 47.095 ;
		RECT	2.58 46.965 2.63 47.095 ;
		RECT	3.84 46.965 3.89 47.095 ;
		RECT	5.675 46.965 5.725 47.095 ;
		RECT	3.06 46.735 3.11 46.865 ;
		RECT	1.085 46.275 1.135 46.405 ;
		RECT	1.405 46.315 1.455 46.365 ;
		RECT	4.47 46.315 4.6 46.365 ;
		RECT	3.06 44.315 3.11 44.445 ;
		RECT	1.57 44.085 1.62 44.215 ;
		RECT	2.58 44.085 2.63 44.215 ;
		RECT	3.84 44.085 3.89 44.215 ;
		RECT	5.675 44.085 5.725 44.215 ;
		RECT	3.06 43.855 3.11 43.985 ;
		RECT	1.085 43.395 1.135 43.525 ;
		RECT	1.405 43.435 1.455 43.485 ;
		RECT	4.47 43.435 4.6 43.485 ;
		RECT	3.06 41.435 3.11 41.565 ;
		RECT	1.57 41.205 1.62 41.335 ;
		RECT	2.58 41.205 2.63 41.335 ;
		RECT	3.84 41.205 3.89 41.335 ;
		RECT	5.675 41.205 5.725 41.335 ;
		RECT	3.06 170.575 3.11 170.705 ;
		RECT	1.085 170.115 1.135 170.245 ;
		RECT	1.405 170.155 1.455 170.205 ;
		RECT	4.47 170.155 4.6 170.205 ;
		RECT	3.06 168.155 3.11 168.285 ;
		RECT	1.57 167.925 1.62 168.055 ;
		RECT	2.58 167.925 2.63 168.055 ;
		RECT	3.84 167.925 3.89 168.055 ;
		RECT	5.675 167.925 5.725 168.055 ;
		RECT	3.06 40.975 3.11 41.105 ;
		RECT	1.085 40.515 1.135 40.645 ;
		RECT	1.405 40.555 1.455 40.605 ;
		RECT	4.47 40.555 4.6 40.605 ;
		RECT	3.06 38.555 3.11 38.685 ;
		RECT	1.57 38.325 1.62 38.455 ;
		RECT	2.58 38.325 2.63 38.455 ;
		RECT	3.84 38.325 3.89 38.455 ;
		RECT	5.675 38.325 5.725 38.455 ;
		RECT	3.06 38.095 3.11 38.225 ;
		RECT	1.085 37.635 1.135 37.765 ;
		RECT	1.405 37.675 1.455 37.725 ;
		RECT	4.47 37.675 4.6 37.725 ;
		RECT	3.06 35.675 3.11 35.805 ;
		RECT	1.57 35.445 1.62 35.575 ;
		RECT	2.58 35.445 2.63 35.575 ;
		RECT	3.84 35.445 3.89 35.575 ;
		RECT	5.675 35.445 5.725 35.575 ;
		RECT	3.06 35.215 3.11 35.345 ;
		RECT	1.085 34.755 1.135 34.885 ;
		RECT	1.405 34.795 1.455 34.845 ;
		RECT	4.47 34.795 4.6 34.845 ;
		RECT	3.06 32.795 3.11 32.925 ;
		RECT	1.57 32.565 1.62 32.695 ;
		RECT	2.58 32.565 2.63 32.695 ;
		RECT	3.84 32.565 3.89 32.695 ;
		RECT	5.675 32.565 5.725 32.695 ;
		RECT	3.06 32.335 3.11 32.465 ;
		RECT	1.085 31.875 1.135 32.005 ;
		RECT	1.405 31.915 1.455 31.965 ;
		RECT	4.47 31.915 4.6 31.965 ;
		RECT	3.06 29.915 3.11 30.045 ;
		RECT	1.57 29.685 1.62 29.815 ;
		RECT	2.58 29.685 2.63 29.815 ;
		RECT	3.84 29.685 3.89 29.815 ;
		RECT	5.675 29.685 5.725 29.815 ;
		RECT	3.06 29.455 3.11 29.585 ;
		RECT	1.085 28.995 1.135 29.125 ;
		RECT	1.405 29.035 1.455 29.085 ;
		RECT	4.47 29.035 4.6 29.085 ;
		RECT	3.06 27.035 3.11 27.165 ;
		RECT	1.57 26.805 1.62 26.935 ;
		RECT	2.58 26.805 2.63 26.935 ;
		RECT	3.84 26.805 3.89 26.935 ;
		RECT	5.675 26.805 5.725 26.935 ;
		RECT	3.06 26.575 3.11 26.705 ;
		RECT	1.085 26.115 1.135 26.245 ;
		RECT	1.405 26.155 1.455 26.205 ;
		RECT	4.47 26.155 4.6 26.205 ;
		RECT	3.06 24.155 3.11 24.285 ;
		RECT	1.57 23.925 1.62 24.055 ;
		RECT	2.58 23.925 2.63 24.055 ;
		RECT	3.84 23.925 3.89 24.055 ;
		RECT	5.675 23.925 5.725 24.055 ;
		RECT	3.06 23.695 3.11 23.825 ;
		RECT	1.085 23.235 1.135 23.365 ;
		RECT	1.405 23.275 1.455 23.325 ;
		RECT	4.47 23.275 4.6 23.325 ;
		RECT	3.06 21.275 3.11 21.405 ;
		RECT	1.57 21.045 1.62 21.175 ;
		RECT	2.58 21.045 2.63 21.175 ;
		RECT	3.84 21.045 3.89 21.175 ;
		RECT	5.675 21.045 5.725 21.175 ;
		RECT	3.06 20.815 3.11 20.945 ;
		RECT	1.085 20.355 1.135 20.485 ;
		RECT	1.405 20.395 1.455 20.445 ;
		RECT	4.47 20.395 4.6 20.445 ;
		RECT	3.06 18.395 3.11 18.525 ;
		RECT	1.57 18.165 1.62 18.295 ;
		RECT	2.58 18.165 2.63 18.295 ;
		RECT	3.84 18.165 3.89 18.295 ;
		RECT	5.675 18.165 5.725 18.295 ;
		RECT	3.06 17.935 3.11 18.065 ;
		RECT	1.085 17.475 1.135 17.605 ;
		RECT	1.405 17.515 1.455 17.565 ;
		RECT	4.47 17.515 4.6 17.565 ;
		RECT	3.06 15.515 3.11 15.645 ;
		RECT	1.57 15.285 1.62 15.415 ;
		RECT	2.58 15.285 2.63 15.415 ;
		RECT	3.84 15.285 3.89 15.415 ;
		RECT	5.675 15.285 5.725 15.415 ;
		RECT	3.06 15.055 3.11 15.185 ;
		RECT	1.085 14.595 1.135 14.725 ;
		RECT	1.405 14.635 1.455 14.685 ;
		RECT	4.47 14.635 4.6 14.685 ;
		RECT	3.06 12.635 3.11 12.765 ;
		RECT	1.57 12.405 1.62 12.535 ;
		RECT	2.58 12.405 2.63 12.535 ;
		RECT	3.84 12.405 3.89 12.535 ;
		RECT	5.675 12.405 5.725 12.535 ;
		RECT	3.06 167.695 3.11 167.825 ;
		RECT	1.085 167.235 1.135 167.365 ;
		RECT	1.405 167.275 1.455 167.325 ;
		RECT	4.47 167.275 4.6 167.325 ;
		RECT	3.06 165.275 3.11 165.405 ;
		RECT	1.57 165.045 1.62 165.175 ;
		RECT	2.58 165.045 2.63 165.175 ;
		RECT	3.84 165.045 3.89 165.175 ;
		RECT	5.675 165.045 5.725 165.175 ;
		RECT	3.06 12.175 3.11 12.305 ;
		RECT	1.085 11.715 1.135 11.845 ;
		RECT	1.405 11.755 1.455 11.805 ;
		RECT	4.47 11.755 4.6 11.805 ;
		RECT	3.06 9.755 3.11 9.885 ;
		RECT	1.57 9.525 1.62 9.655 ;
		RECT	2.58 9.525 2.63 9.655 ;
		RECT	3.84 9.525 3.89 9.655 ;
		RECT	5.675 9.525 5.725 9.655 ;
		RECT	3.06 9.295 3.11 9.425 ;
		RECT	1.085 8.835 1.135 8.965 ;
		RECT	1.405 8.875 1.455 8.925 ;
		RECT	4.47 8.875 4.6 8.925 ;
		RECT	3.06 6.875 3.11 7.005 ;
		RECT	1.57 6.645 1.62 6.775 ;
		RECT	2.58 6.645 2.63 6.775 ;
		RECT	3.84 6.645 3.89 6.775 ;
		RECT	5.675 6.645 5.725 6.775 ;
		RECT	3.06 6.415 3.11 6.545 ;
		RECT	1.085 5.955 1.135 6.085 ;
		RECT	1.405 5.995 1.455 6.045 ;
		RECT	4.47 5.995 4.6 6.045 ;
		RECT	3.06 3.995 3.11 4.125 ;
		RECT	1.57 3.765 1.62 3.895 ;
		RECT	2.58 3.765 2.63 3.895 ;
		RECT	3.84 3.765 3.89 3.895 ;
		RECT	5.675 3.765 5.725 3.895 ;
		RECT	3.06 164.815 3.11 164.945 ;
		RECT	1.085 164.355 1.135 164.485 ;
		RECT	1.405 164.395 1.455 164.445 ;
		RECT	4.47 164.395 4.6 164.445 ;
		RECT	3.06 162.395 3.11 162.525 ;
		RECT	1.57 162.165 1.62 162.295 ;
		RECT	2.58 162.165 2.63 162.295 ;
		RECT	3.84 162.165 3.89 162.295 ;
		RECT	5.675 162.165 5.725 162.295 ;
		RECT	3.06 161.935 3.11 162.065 ;
		RECT	1.085 161.475 1.135 161.605 ;
		RECT	1.405 161.515 1.455 161.565 ;
		RECT	4.47 161.515 4.6 161.565 ;
		RECT	3.06 159.515 3.11 159.645 ;
		RECT	1.57 159.285 1.62 159.415 ;
		RECT	2.58 159.285 2.63 159.415 ;
		RECT	3.84 159.285 3.89 159.415 ;
		RECT	5.675 159.285 5.725 159.415 ;
		RECT	3.06 159.055 3.11 159.185 ;
		RECT	1.085 158.595 1.135 158.725 ;
		RECT	1.405 158.635 1.455 158.685 ;
		RECT	4.47 158.635 4.6 158.685 ;
		RECT	3.06 156.635 3.11 156.765 ;
		RECT	1.57 156.405 1.62 156.535 ;
		RECT	2.58 156.405 2.63 156.535 ;
		RECT	3.84 156.405 3.89 156.535 ;
		RECT	5.675 156.405 5.725 156.535 ;
		RECT	3.06 3.535 3.11 3.665 ;
		RECT	1.085 3.075 1.135 3.205 ;
		RECT	1.405 3.115 1.455 3.165 ;
		RECT	4.47 3.115 4.6 3.165 ;
		RECT	3.06 1.115 3.11 1.245 ;
		RECT	1.57 0.885 1.62 1.015 ;
		RECT	2.58 0.885 2.63 1.015 ;
		RECT	3.84 0.885 3.89 1.015 ;
		RECT	5.675 0.885 5.725 1.015 ;
		RECT	3.06 184.975 3.11 185.105 ;
		RECT	1.085 184.515 1.135 184.645 ;
		RECT	1.405 184.555 1.455 184.605 ;
		RECT	4.47 184.555 4.6 184.605 ;
		RECT	3.06 182.555 3.11 182.685 ;
		RECT	1.57 182.325 1.62 182.455 ;
		RECT	2.58 182.325 2.63 182.455 ;
		RECT	3.84 182.325 3.89 182.455 ;
		RECT	5.675 182.325 5.725 182.455 ;
		RECT	0.435 184.515 0.485 184.645 ;
		RECT	0.435 184.975 0.485 185.105 ;
		RECT	0.435 182.555 0.485 182.685 ;
		RECT	0.435 181.635 0.485 181.765 ;
		RECT	0.435 182.095 0.485 182.225 ;
		RECT	0.435 179.675 0.485 179.805 ;
		RECT	0.435 155.715 0.485 155.845 ;
		RECT	0.435 156.175 0.485 156.305 ;
		RECT	0.435 153.755 0.485 153.885 ;
		RECT	0.435 152.835 0.485 152.965 ;
		RECT	0.435 153.295 0.485 153.425 ;
		RECT	0.435 150.875 0.485 151.005 ;
		RECT	0.435 149.955 0.485 150.085 ;
		RECT	0.435 150.415 0.485 150.545 ;
		RECT	0.435 147.995 0.485 148.125 ;
		RECT	0.435 147.075 0.485 147.205 ;
		RECT	0.435 147.535 0.485 147.665 ;
		RECT	0.435 145.115 0.485 145.245 ;
		RECT	0.435 144.195 0.485 144.325 ;
		RECT	0.435 144.655 0.485 144.785 ;
		RECT	0.435 142.235 0.485 142.365 ;
		RECT	0.435 141.315 0.485 141.445 ;
		RECT	0.435 141.775 0.485 141.905 ;
		RECT	0.435 139.355 0.485 139.485 ;
		RECT	0.435 138.435 0.485 138.565 ;
		RECT	0.435 138.895 0.485 139.025 ;
		RECT	0.435 136.475 0.485 136.605 ;
		RECT	0.435 135.555 0.485 135.685 ;
		RECT	0.435 136.015 0.485 136.145 ;
		RECT	0.435 133.595 0.485 133.725 ;
		RECT	0.435 132.675 0.485 132.805 ;
		RECT	0.435 133.135 0.485 133.265 ;
		RECT	0.435 130.715 0.485 130.845 ;
		RECT	0.435 129.795 0.485 129.925 ;
		RECT	0.435 130.255 0.485 130.385 ;
		RECT	0.435 127.835 0.485 127.965 ;
		RECT	0.435 178.755 0.485 178.885 ;
		RECT	0.435 179.215 0.485 179.345 ;
		RECT	0.435 176.795 0.485 176.925 ;
		RECT	0.435 126.915 0.485 127.045 ;
		RECT	0.435 127.375 0.485 127.505 ;
		RECT	0.435 124.955 0.485 125.085 ;
		RECT	0.435 124.035 0.485 124.165 ;
		RECT	0.435 124.495 0.485 124.625 ;
		RECT	0.435 122.075 0.485 122.205 ;
		RECT	0.435 121.155 0.485 121.285 ;
		RECT	0.435 121.615 0.485 121.745 ;
		RECT	0.435 119.195 0.485 119.325 ;
		RECT	0.435 118.275 0.485 118.405 ;
		RECT	0.435 118.735 0.485 118.865 ;
		RECT	0.435 116.315 0.485 116.445 ;
		RECT	0.435 115.395 0.485 115.525 ;
		RECT	0.435 115.855 0.485 115.985 ;
		RECT	0.435 113.435 0.485 113.565 ;
		RECT	0.435 112.515 0.485 112.645 ;
		RECT	0.435 112.975 0.485 113.105 ;
		RECT	0.435 110.555 0.485 110.685 ;
		RECT	0.435 109.635 0.485 109.765 ;
		RECT	0.435 110.095 0.485 110.225 ;
		RECT	0.435 107.675 0.485 107.805 ;
		RECT	0.435 106.755 0.485 106.885 ;
		RECT	0.435 107.215 0.485 107.345 ;
		RECT	0.435 104.795 0.485 104.925 ;
		RECT	0.435 103.875 0.485 104.005 ;
		RECT	0.435 104.335 0.485 104.465 ;
		RECT	0.435 101.915 0.485 102.045 ;
		RECT	0.435 100.995 0.485 101.125 ;
		RECT	0.435 101.455 0.485 101.585 ;
		RECT	0.435 99.035 0.485 99.165 ;
		RECT	0.435 175.875 0.485 176.005 ;
		RECT	0.435 176.335 0.485 176.465 ;
		RECT	0.435 173.915 0.485 174.045 ;
		RECT	0.435 98.115 0.485 98.245 ;
		RECT	0.435 98.575 0.485 98.705 ;
		RECT	0.435 96.155 0.485 96.285 ;
		RECT	0.435 95.235 0.485 95.365 ;
		RECT	0.435 95.695 0.485 95.825 ;
		RECT	0.435 93.275 0.485 93.405 ;
		RECT	0.435 92.355 0.485 92.485 ;
		RECT	0.435 92.815 0.485 92.945 ;
		RECT	0.435 90.395 0.485 90.525 ;
		RECT	0.435 89.475 0.485 89.605 ;
		RECT	0.435 89.935 0.485 90.065 ;
		RECT	0.435 87.515 0.485 87.645 ;
		RECT	0.435 86.595 0.485 86.725 ;
		RECT	0.435 87.055 0.485 87.185 ;
		RECT	0.435 84.635 0.485 84.765 ;
		RECT	0.435 83.715 0.485 83.845 ;
		RECT	0.435 84.175 0.485 84.305 ;
		RECT	0.435 81.755 0.485 81.885 ;
		RECT	0.435 80.835 0.485 80.965 ;
		RECT	0.435 81.295 0.485 81.425 ;
		RECT	0.435 78.875 0.485 79.005 ;
		RECT	0.435 77.955 0.485 78.085 ;
		RECT	0.435 78.415 0.485 78.545 ;
		RECT	0.435 75.995 0.485 76.125 ;
		RECT	0.435 75.075 0.485 75.205 ;
		RECT	0.435 75.535 0.485 75.665 ;
		RECT	0.435 73.115 0.485 73.245 ;
		RECT	0.435 72.195 0.485 72.325 ;
		RECT	0.435 72.655 0.485 72.785 ;
		RECT	0.435 70.235 0.485 70.365 ;
		RECT	0.435 172.995 0.485 173.125 ;
		RECT	0.435 173.455 0.485 173.585 ;
		RECT	0.435 171.035 0.485 171.165 ;
		RECT	0.435 69.315 0.485 69.445 ;
		RECT	0.435 69.775 0.485 69.905 ;
		RECT	0.435 67.355 0.485 67.485 ;
		RECT	0.435 66.435 0.485 66.565 ;
		RECT	0.435 66.895 0.485 67.025 ;
		RECT	0.435 64.475 0.485 64.605 ;
		RECT	0.435 63.555 0.485 63.685 ;
		RECT	0.435 64.015 0.485 64.145 ;
		RECT	0.435 61.595 0.485 61.725 ;
		RECT	0.435 60.675 0.485 60.805 ;
		RECT	0.435 61.135 0.485 61.265 ;
		RECT	0.435 58.715 0.485 58.845 ;
		RECT	0.435 57.795 0.485 57.925 ;
		RECT	0.435 58.255 0.485 58.385 ;
		RECT	0.435 55.835 0.485 55.965 ;
		RECT	0.435 54.915 0.485 55.045 ;
		RECT	0.435 55.375 0.485 55.505 ;
		RECT	0.435 52.955 0.485 53.085 ;
		RECT	0.435 52.035 0.485 52.165 ;
		RECT	0.435 52.495 0.485 52.625 ;
		RECT	0.435 50.075 0.485 50.205 ;
		RECT	0.435 49.155 0.485 49.285 ;
		RECT	0.435 49.615 0.485 49.745 ;
		RECT	0.435 47.195 0.485 47.325 ;
		RECT	0.435 46.275 0.485 46.405 ;
		RECT	0.435 46.735 0.485 46.865 ;
		RECT	0.435 44.315 0.485 44.445 ;
		RECT	0.435 43.395 0.485 43.525 ;
		RECT	0.435 43.855 0.485 43.985 ;
		RECT	0.435 41.435 0.485 41.565 ;
		RECT	0.435 170.115 0.485 170.245 ;
		RECT	0.435 170.575 0.485 170.705 ;
		RECT	0.435 168.155 0.485 168.285 ;
		RECT	0.435 40.515 0.485 40.645 ;
		RECT	0.435 40.975 0.485 41.105 ;
		RECT	0.435 38.555 0.485 38.685 ;
		RECT	0.435 37.635 0.485 37.765 ;
		RECT	0.435 38.095 0.485 38.225 ;
		RECT	0.435 35.675 0.485 35.805 ;
		RECT	0.435 34.755 0.485 34.885 ;
		RECT	0.435 35.215 0.485 35.345 ;
		RECT	0.435 32.795 0.485 32.925 ;
		RECT	0.435 31.875 0.485 32.005 ;
		RECT	0.435 32.335 0.485 32.465 ;
		RECT	0.435 29.915 0.485 30.045 ;
		RECT	0.435 28.995 0.485 29.125 ;
		RECT	0.435 29.455 0.485 29.585 ;
		RECT	0.435 27.035 0.485 27.165 ;
		RECT	0.435 26.115 0.485 26.245 ;
		RECT	0.435 26.575 0.485 26.705 ;
		RECT	0.435 24.155 0.485 24.285 ;
		RECT	0.435 23.235 0.485 23.365 ;
		RECT	0.435 23.695 0.485 23.825 ;
		RECT	0.435 21.275 0.485 21.405 ;
		RECT	0.435 20.355 0.485 20.485 ;
		RECT	0.435 20.815 0.485 20.945 ;
		RECT	0.435 18.395 0.485 18.525 ;
		RECT	0.435 17.475 0.485 17.605 ;
		RECT	0.435 17.935 0.485 18.065 ;
		RECT	0.435 15.515 0.485 15.645 ;
		RECT	0.435 14.595 0.485 14.725 ;
		RECT	0.435 15.055 0.485 15.185 ;
		RECT	0.435 12.635 0.485 12.765 ;
		RECT	0.435 167.235 0.485 167.365 ;
		RECT	0.435 167.695 0.485 167.825 ;
		RECT	0.435 165.275 0.485 165.405 ;
		RECT	0.435 11.715 0.485 11.845 ;
		RECT	0.435 12.175 0.485 12.305 ;
		RECT	0.435 9.755 0.485 9.885 ;
		RECT	0.435 8.835 0.485 8.965 ;
		RECT	0.435 9.295 0.485 9.425 ;
		RECT	0.435 6.875 0.485 7.005 ;
		RECT	0.435 5.955 0.485 6.085 ;
		RECT	0.435 6.415 0.485 6.545 ;
		RECT	0.435 3.995 0.485 4.125 ;
		RECT	0.435 3.075 0.485 3.205 ;
		RECT	0.435 3.535 0.485 3.665 ;
		RECT	0.435 1.115 0.485 1.245 ;
		RECT	0.435 164.355 0.485 164.485 ;
		RECT	0.435 164.815 0.485 164.945 ;
		RECT	0.435 162.395 0.485 162.525 ;
		RECT	0.435 161.475 0.485 161.605 ;
		RECT	0.435 161.935 0.485 162.065 ;
		RECT	0.435 159.515 0.485 159.645 ;
		RECT	0.435 158.595 0.485 158.725 ;
		RECT	0.435 159.055 0.485 159.185 ;
		RECT	0.435 156.635 0.485 156.765 ;
		RECT	6.22 229.755 6.27 229.885 ;
		RECT	7.5 229.755 7.55 229.885 ;
		RECT	9.04 229.755 9.09 229.885 ;
		RECT	9.315 229.755 9.365 229.885 ;
		RECT	9.72 229.755 9.77 229.885 ;
		RECT	11.025 229.755 11.075 229.885 ;
		RECT	12.79 229.755 12.84 229.885 ;
		RECT	6.225 232.175 6.275 232.305 ;
		RECT	7.5 232.175 7.55 232.305 ;
		RECT	9.04 232.175 9.09 232.305 ;
		RECT	9.315 232.175 9.365 232.305 ;
		RECT	11.025 232.175 11.075 232.305 ;
		RECT	12.79 232.175 12.84 232.305 ;
		RECT	7.18 232.405 7.23 232.535 ;
		RECT	14.14 232.405 14.19 232.535 ;
		RECT	8.56 229.755 8.61 229.885 ;
		RECT	10.27 229.755 10.32 229.885 ;
		RECT	8.56 232.175 8.61 232.305 ;
		RECT	10.27 232.175 10.32 232.305 ;
		RECT	6.22 232.635 6.27 232.765 ;
		RECT	7.5 232.635 7.55 232.765 ;
		RECT	9.04 232.635 9.09 232.765 ;
		RECT	9.315 232.635 9.365 232.765 ;
		RECT	9.72 232.635 9.77 232.765 ;
		RECT	11.025 232.635 11.075 232.765 ;
		RECT	12.79 232.635 12.84 232.765 ;
		RECT	6.225 235.055 6.275 235.185 ;
		RECT	7.5 235.055 7.55 235.185 ;
		RECT	9.04 235.055 9.09 235.185 ;
		RECT	9.315 235.055 9.365 235.185 ;
		RECT	11.025 235.055 11.075 235.185 ;
		RECT	12.79 235.055 12.84 235.185 ;
		RECT	7.18 235.285 7.23 235.415 ;
		RECT	14.14 235.285 14.19 235.415 ;
		RECT	8.56 232.635 8.61 232.765 ;
		RECT	10.27 232.635 10.32 232.765 ;
		RECT	8.56 235.055 8.61 235.185 ;
		RECT	10.27 235.055 10.32 235.185 ;
		RECT	6.22 235.515 6.27 235.645 ;
		RECT	7.5 235.515 7.55 235.645 ;
		RECT	9.04 235.515 9.09 235.645 ;
		RECT	9.315 235.515 9.365 235.645 ;
		RECT	9.72 235.515 9.77 235.645 ;
		RECT	11.025 235.515 11.075 235.645 ;
		RECT	12.79 235.515 12.84 235.645 ;
		RECT	6.225 237.935 6.275 238.065 ;
		RECT	7.5 237.935 7.55 238.065 ;
		RECT	9.04 237.935 9.09 238.065 ;
		RECT	9.315 237.935 9.365 238.065 ;
		RECT	11.025 237.935 11.075 238.065 ;
		RECT	12.79 237.935 12.84 238.065 ;
		RECT	7.18 238.165 7.23 238.295 ;
		RECT	14.14 238.165 14.19 238.295 ;
		RECT	8.56 235.515 8.61 235.645 ;
		RECT	10.27 235.515 10.32 235.645 ;
		RECT	8.56 237.935 8.61 238.065 ;
		RECT	10.27 237.935 10.32 238.065 ;
		RECT	6.22 238.395 6.27 238.525 ;
		RECT	7.5 238.395 7.55 238.525 ;
		RECT	9.04 238.395 9.09 238.525 ;
		RECT	9.315 238.395 9.365 238.525 ;
		RECT	9.72 238.395 9.77 238.525 ;
		RECT	11.025 238.395 11.075 238.525 ;
		RECT	12.79 238.395 12.84 238.525 ;
		RECT	6.225 240.815 6.275 240.945 ;
		RECT	7.5 240.815 7.55 240.945 ;
		RECT	9.04 240.815 9.09 240.945 ;
		RECT	9.315 240.815 9.365 240.945 ;
		RECT	11.025 240.815 11.075 240.945 ;
		RECT	12.79 240.815 12.84 240.945 ;
		RECT	7.18 241.045 7.23 241.175 ;
		RECT	14.14 241.045 14.19 241.175 ;
		RECT	8.56 238.395 8.61 238.525 ;
		RECT	10.27 238.395 10.32 238.525 ;
		RECT	8.56 240.815 8.61 240.945 ;
		RECT	10.27 240.815 10.32 240.945 ;
		RECT	6.22 241.275 6.27 241.405 ;
		RECT	7.5 241.275 7.55 241.405 ;
		RECT	9.04 241.275 9.09 241.405 ;
		RECT	9.315 241.275 9.365 241.405 ;
		RECT	9.72 241.275 9.77 241.405 ;
		RECT	11.025 241.275 11.075 241.405 ;
		RECT	12.79 241.275 12.84 241.405 ;
		RECT	6.225 243.695 6.275 243.825 ;
		RECT	7.5 243.695 7.55 243.825 ;
		RECT	9.04 243.695 9.09 243.825 ;
		RECT	9.315 243.695 9.365 243.825 ;
		RECT	11.025 243.695 11.075 243.825 ;
		RECT	12.79 243.695 12.84 243.825 ;
		RECT	7.18 243.925 7.23 244.055 ;
		RECT	14.14 243.925 14.19 244.055 ;
		RECT	8.56 241.275 8.61 241.405 ;
		RECT	10.27 241.275 10.32 241.405 ;
		RECT	8.56 243.695 8.61 243.825 ;
		RECT	10.27 243.695 10.32 243.825 ;
		RECT	6.22 244.155 6.27 244.285 ;
		RECT	7.5 244.155 7.55 244.285 ;
		RECT	9.04 244.155 9.09 244.285 ;
		RECT	9.315 244.155 9.365 244.285 ;
		RECT	9.72 244.155 9.77 244.285 ;
		RECT	11.025 244.155 11.075 244.285 ;
		RECT	12.79 244.155 12.84 244.285 ;
		RECT	6.225 246.575 6.275 246.705 ;
		RECT	7.5 246.575 7.55 246.705 ;
		RECT	9.04 246.575 9.09 246.705 ;
		RECT	9.315 246.575 9.365 246.705 ;
		RECT	11.025 246.575 11.075 246.705 ;
		RECT	12.79 246.575 12.84 246.705 ;
		RECT	7.18 246.805 7.23 246.935 ;
		RECT	14.14 246.805 14.19 246.935 ;
		RECT	8.56 244.155 8.61 244.285 ;
		RECT	10.27 244.155 10.32 244.285 ;
		RECT	8.56 246.575 8.61 246.705 ;
		RECT	10.27 246.575 10.32 246.705 ;
		RECT	6.22 247.035 6.27 247.165 ;
		RECT	7.5 247.035 7.55 247.165 ;
		RECT	9.04 247.035 9.09 247.165 ;
		RECT	9.315 247.035 9.365 247.165 ;
		RECT	9.72 247.035 9.77 247.165 ;
		RECT	11.025 247.035 11.075 247.165 ;
		RECT	12.79 247.035 12.84 247.165 ;
		RECT	6.225 249.455 6.275 249.585 ;
		RECT	7.5 249.455 7.55 249.585 ;
		RECT	9.04 249.455 9.09 249.585 ;
		RECT	9.315 249.455 9.365 249.585 ;
		RECT	11.025 249.455 11.075 249.585 ;
		RECT	12.79 249.455 12.84 249.585 ;
		RECT	7.18 249.685 7.23 249.815 ;
		RECT	14.14 249.685 14.19 249.815 ;
		RECT	8.56 247.035 8.61 247.165 ;
		RECT	10.27 247.035 10.32 247.165 ;
		RECT	8.56 249.455 8.61 249.585 ;
		RECT	10.27 249.455 10.32 249.585 ;
		RECT	6.22 249.915 6.27 250.045 ;
		RECT	7.5 249.915 7.55 250.045 ;
		RECT	9.04 249.915 9.09 250.045 ;
		RECT	9.315 249.915 9.365 250.045 ;
		RECT	9.72 249.915 9.77 250.045 ;
		RECT	11.025 249.915 11.075 250.045 ;
		RECT	12.79 249.915 12.84 250.045 ;
		RECT	6.225 252.335 6.275 252.465 ;
		RECT	7.5 252.335 7.55 252.465 ;
		RECT	9.04 252.335 9.09 252.465 ;
		RECT	9.315 252.335 9.365 252.465 ;
		RECT	11.025 252.335 11.075 252.465 ;
		RECT	12.79 252.335 12.84 252.465 ;
		RECT	7.18 252.565 7.23 252.695 ;
		RECT	14.14 252.565 14.19 252.695 ;
		RECT	8.56 249.915 8.61 250.045 ;
		RECT	10.27 249.915 10.32 250.045 ;
		RECT	8.56 252.335 8.61 252.465 ;
		RECT	10.27 252.335 10.32 252.465 ;
		RECT	6.22 252.795 6.27 252.925 ;
		RECT	7.5 252.795 7.55 252.925 ;
		RECT	9.04 252.795 9.09 252.925 ;
		RECT	9.315 252.795 9.365 252.925 ;
		RECT	9.72 252.795 9.77 252.925 ;
		RECT	11.025 252.795 11.075 252.925 ;
		RECT	12.79 252.795 12.84 252.925 ;
		RECT	6.225 255.215 6.275 255.345 ;
		RECT	7.5 255.215 7.55 255.345 ;
		RECT	9.04 255.215 9.09 255.345 ;
		RECT	9.315 255.215 9.365 255.345 ;
		RECT	11.025 255.215 11.075 255.345 ;
		RECT	12.79 255.215 12.84 255.345 ;
		RECT	7.18 255.445 7.23 255.575 ;
		RECT	14.14 255.445 14.19 255.575 ;
		RECT	8.56 252.795 8.61 252.925 ;
		RECT	10.27 252.795 10.32 252.925 ;
		RECT	8.56 255.215 8.61 255.345 ;
		RECT	10.27 255.215 10.32 255.345 ;
		RECT	6.22 255.675 6.27 255.805 ;
		RECT	7.5 255.675 7.55 255.805 ;
		RECT	9.04 255.675 9.09 255.805 ;
		RECT	9.315 255.675 9.365 255.805 ;
		RECT	9.72 255.675 9.77 255.805 ;
		RECT	11.025 255.675 11.075 255.805 ;
		RECT	12.79 255.675 12.84 255.805 ;
		RECT	6.225 258.095 6.275 258.225 ;
		RECT	7.5 258.095 7.55 258.225 ;
		RECT	9.04 258.095 9.09 258.225 ;
		RECT	9.315 258.095 9.365 258.225 ;
		RECT	11.025 258.095 11.075 258.225 ;
		RECT	12.79 258.095 12.84 258.225 ;
		RECT	7.18 258.325 7.23 258.455 ;
		RECT	14.14 258.325 14.19 258.455 ;
		RECT	8.56 255.675 8.61 255.805 ;
		RECT	10.27 255.675 10.32 255.805 ;
		RECT	8.56 258.095 8.61 258.225 ;
		RECT	10.27 258.095 10.32 258.225 ;
		RECT	6.22 258.555 6.27 258.685 ;
		RECT	7.5 258.555 7.55 258.685 ;
		RECT	9.04 258.555 9.09 258.685 ;
		RECT	9.315 258.555 9.365 258.685 ;
		RECT	9.72 258.555 9.77 258.685 ;
		RECT	11.025 258.555 11.075 258.685 ;
		RECT	12.79 258.555 12.84 258.685 ;
		RECT	6.225 260.975 6.275 261.105 ;
		RECT	7.5 260.975 7.55 261.105 ;
		RECT	9.04 260.975 9.09 261.105 ;
		RECT	9.315 260.975 9.365 261.105 ;
		RECT	11.025 260.975 11.075 261.105 ;
		RECT	12.79 260.975 12.84 261.105 ;
		RECT	7.18 261.205 7.23 261.335 ;
		RECT	14.14 261.205 14.19 261.335 ;
		RECT	8.56 258.555 8.61 258.685 ;
		RECT	10.27 258.555 10.32 258.685 ;
		RECT	8.56 260.975 8.61 261.105 ;
		RECT	10.27 260.975 10.32 261.105 ;
		RECT	6.22 261.435 6.27 261.565 ;
		RECT	7.5 261.435 7.55 261.565 ;
		RECT	9.04 261.435 9.09 261.565 ;
		RECT	9.315 261.435 9.365 261.565 ;
		RECT	9.72 261.435 9.77 261.565 ;
		RECT	11.025 261.435 11.075 261.565 ;
		RECT	12.79 261.435 12.84 261.565 ;
		RECT	6.225 263.855 6.275 263.985 ;
		RECT	7.5 263.855 7.55 263.985 ;
		RECT	9.04 263.855 9.09 263.985 ;
		RECT	9.315 263.855 9.365 263.985 ;
		RECT	11.025 263.855 11.075 263.985 ;
		RECT	12.79 263.855 12.84 263.985 ;
		RECT	7.18 264.085 7.23 264.215 ;
		RECT	14.14 264.085 14.19 264.215 ;
		RECT	8.56 261.435 8.61 261.565 ;
		RECT	10.27 261.435 10.32 261.565 ;
		RECT	8.56 263.855 8.61 263.985 ;
		RECT	10.27 263.855 10.32 263.985 ;
		RECT	6.22 264.315 6.27 264.445 ;
		RECT	7.5 264.315 7.55 264.445 ;
		RECT	9.04 264.315 9.09 264.445 ;
		RECT	9.315 264.315 9.365 264.445 ;
		RECT	9.72 264.315 9.77 264.445 ;
		RECT	11.025 264.315 11.075 264.445 ;
		RECT	12.79 264.315 12.84 264.445 ;
		RECT	6.225 266.735 6.275 266.865 ;
		RECT	7.5 266.735 7.55 266.865 ;
		RECT	9.04 266.735 9.09 266.865 ;
		RECT	9.315 266.735 9.365 266.865 ;
		RECT	11.025 266.735 11.075 266.865 ;
		RECT	12.79 266.735 12.84 266.865 ;
		RECT	7.18 266.965 7.23 267.095 ;
		RECT	14.14 266.965 14.19 267.095 ;
		RECT	8.56 264.315 8.61 264.445 ;
		RECT	10.27 264.315 10.32 264.445 ;
		RECT	8.56 266.735 8.61 266.865 ;
		RECT	10.27 266.735 10.32 266.865 ;
		RECT	6.22 267.195 6.27 267.325 ;
		RECT	7.5 267.195 7.55 267.325 ;
		RECT	9.04 267.195 9.09 267.325 ;
		RECT	9.315 267.195 9.365 267.325 ;
		RECT	9.72 267.195 9.77 267.325 ;
		RECT	11.025 267.195 11.075 267.325 ;
		RECT	12.79 267.195 12.84 267.325 ;
		RECT	6.225 269.615 6.275 269.745 ;
		RECT	7.5 269.615 7.55 269.745 ;
		RECT	9.04 269.615 9.09 269.745 ;
		RECT	9.315 269.615 9.365 269.745 ;
		RECT	11.025 269.615 11.075 269.745 ;
		RECT	12.79 269.615 12.84 269.745 ;
		RECT	7.18 269.845 7.23 269.975 ;
		RECT	14.14 269.845 14.19 269.975 ;
		RECT	8.56 267.195 8.61 267.325 ;
		RECT	10.27 267.195 10.32 267.325 ;
		RECT	8.56 269.615 8.61 269.745 ;
		RECT	10.27 269.615 10.32 269.745 ;
		RECT	6.22 270.075 6.27 270.205 ;
		RECT	7.5 270.075 7.55 270.205 ;
		RECT	9.04 270.075 9.09 270.205 ;
		RECT	9.315 270.075 9.365 270.205 ;
		RECT	9.72 270.075 9.77 270.205 ;
		RECT	11.025 270.075 11.075 270.205 ;
		RECT	12.79 270.075 12.84 270.205 ;
		RECT	6.225 272.495 6.275 272.625 ;
		RECT	7.5 272.495 7.55 272.625 ;
		RECT	9.04 272.495 9.09 272.625 ;
		RECT	9.315 272.495 9.365 272.625 ;
		RECT	11.025 272.495 11.075 272.625 ;
		RECT	12.79 272.495 12.84 272.625 ;
		RECT	7.18 272.725 7.23 272.855 ;
		RECT	14.14 272.725 14.19 272.855 ;
		RECT	8.56 270.075 8.61 270.205 ;
		RECT	10.27 270.075 10.32 270.205 ;
		RECT	8.56 272.495 8.61 272.625 ;
		RECT	10.27 272.495 10.32 272.625 ;
		RECT	6.22 272.955 6.27 273.085 ;
		RECT	7.5 272.955 7.55 273.085 ;
		RECT	9.04 272.955 9.09 273.085 ;
		RECT	9.315 272.955 9.365 273.085 ;
		RECT	9.72 272.955 9.77 273.085 ;
		RECT	11.025 272.955 11.075 273.085 ;
		RECT	12.79 272.955 12.84 273.085 ;
		RECT	6.225 275.375 6.275 275.505 ;
		RECT	7.5 275.375 7.55 275.505 ;
		RECT	9.04 275.375 9.09 275.505 ;
		RECT	9.315 275.375 9.365 275.505 ;
		RECT	11.025 275.375 11.075 275.505 ;
		RECT	12.79 275.375 12.84 275.505 ;
		RECT	7.18 275.605 7.23 275.735 ;
		RECT	14.14 275.605 14.19 275.735 ;
		RECT	8.56 272.955 8.61 273.085 ;
		RECT	10.27 272.955 10.32 273.085 ;
		RECT	8.56 275.375 8.61 275.505 ;
		RECT	10.27 275.375 10.32 275.505 ;
		RECT	6.22 275.835 6.27 275.965 ;
		RECT	7.5 275.835 7.55 275.965 ;
		RECT	9.04 275.835 9.09 275.965 ;
		RECT	9.315 275.835 9.365 275.965 ;
		RECT	9.72 275.835 9.77 275.965 ;
		RECT	11.025 275.835 11.075 275.965 ;
		RECT	12.79 275.835 12.84 275.965 ;
		RECT	6.225 278.255 6.275 278.385 ;
		RECT	7.5 278.255 7.55 278.385 ;
		RECT	9.04 278.255 9.09 278.385 ;
		RECT	9.315 278.255 9.365 278.385 ;
		RECT	11.025 278.255 11.075 278.385 ;
		RECT	12.79 278.255 12.84 278.385 ;
		RECT	7.18 278.485 7.23 278.615 ;
		RECT	14.14 278.485 14.19 278.615 ;
		RECT	8.56 275.835 8.61 275.965 ;
		RECT	10.27 275.835 10.32 275.965 ;
		RECT	8.56 278.255 8.61 278.385 ;
		RECT	10.27 278.255 10.32 278.385 ;
		RECT	6.22 278.715 6.27 278.845 ;
		RECT	7.5 278.715 7.55 278.845 ;
		RECT	9.04 278.715 9.09 278.845 ;
		RECT	9.315 278.715 9.365 278.845 ;
		RECT	9.72 278.715 9.77 278.845 ;
		RECT	11.025 278.715 11.075 278.845 ;
		RECT	12.79 278.715 12.84 278.845 ;
		RECT	6.225 281.135 6.275 281.265 ;
		RECT	7.5 281.135 7.55 281.265 ;
		RECT	9.04 281.135 9.09 281.265 ;
		RECT	9.315 281.135 9.365 281.265 ;
		RECT	11.025 281.135 11.075 281.265 ;
		RECT	12.79 281.135 12.84 281.265 ;
		RECT	7.18 281.365 7.23 281.495 ;
		RECT	14.14 281.365 14.19 281.495 ;
		RECT	8.56 278.715 8.61 278.845 ;
		RECT	10.27 278.715 10.32 278.845 ;
		RECT	8.56 281.135 8.61 281.265 ;
		RECT	10.27 281.135 10.32 281.265 ;
		RECT	6.22 281.595 6.27 281.725 ;
		RECT	7.5 281.595 7.55 281.725 ;
		RECT	9.04 281.595 9.09 281.725 ;
		RECT	9.315 281.595 9.365 281.725 ;
		RECT	9.72 281.595 9.77 281.725 ;
		RECT	11.025 281.595 11.075 281.725 ;
		RECT	12.79 281.595 12.84 281.725 ;
		RECT	6.225 284.015 6.275 284.145 ;
		RECT	7.5 284.015 7.55 284.145 ;
		RECT	9.04 284.015 9.09 284.145 ;
		RECT	9.315 284.015 9.365 284.145 ;
		RECT	11.025 284.015 11.075 284.145 ;
		RECT	12.79 284.015 12.84 284.145 ;
		RECT	7.18 284.245 7.23 284.375 ;
		RECT	14.14 284.245 14.19 284.375 ;
		RECT	8.56 281.595 8.61 281.725 ;
		RECT	10.27 281.595 10.32 281.725 ;
		RECT	8.56 284.015 8.61 284.145 ;
		RECT	10.27 284.015 10.32 284.145 ;
		RECT	6.22 284.475 6.27 284.605 ;
		RECT	7.5 284.475 7.55 284.605 ;
		RECT	9.04 284.475 9.09 284.605 ;
		RECT	9.315 284.475 9.365 284.605 ;
		RECT	9.72 284.475 9.77 284.605 ;
		RECT	11.025 284.475 11.075 284.605 ;
		RECT	12.79 284.475 12.84 284.605 ;
		RECT	6.225 286.895 6.275 287.025 ;
		RECT	7.5 286.895 7.55 287.025 ;
		RECT	9.04 286.895 9.09 287.025 ;
		RECT	9.315 286.895 9.365 287.025 ;
		RECT	11.025 286.895 11.075 287.025 ;
		RECT	12.79 286.895 12.84 287.025 ;
		RECT	7.18 287.125 7.23 287.255 ;
		RECT	14.14 287.125 14.19 287.255 ;
		RECT	8.56 284.475 8.61 284.605 ;
		RECT	10.27 284.475 10.32 284.605 ;
		RECT	8.56 286.895 8.61 287.025 ;
		RECT	10.27 286.895 10.32 287.025 ;
		RECT	6.22 287.355 6.27 287.485 ;
		RECT	7.5 287.355 7.55 287.485 ;
		RECT	9.04 287.355 9.09 287.485 ;
		RECT	9.315 287.355 9.365 287.485 ;
		RECT	9.72 287.355 9.77 287.485 ;
		RECT	11.025 287.355 11.075 287.485 ;
		RECT	12.79 287.355 12.84 287.485 ;
		RECT	6.225 289.775 6.275 289.905 ;
		RECT	7.5 289.775 7.55 289.905 ;
		RECT	9.04 289.775 9.09 289.905 ;
		RECT	9.315 289.775 9.365 289.905 ;
		RECT	11.025 289.775 11.075 289.905 ;
		RECT	12.79 289.775 12.84 289.905 ;
		RECT	7.18 290.005 7.23 290.135 ;
		RECT	14.14 290.005 14.19 290.135 ;
		RECT	8.56 287.355 8.61 287.485 ;
		RECT	10.27 287.355 10.32 287.485 ;
		RECT	8.56 289.775 8.61 289.905 ;
		RECT	10.27 289.775 10.32 289.905 ;
		RECT	6.22 290.235 6.27 290.365 ;
		RECT	7.5 290.235 7.55 290.365 ;
		RECT	9.04 290.235 9.09 290.365 ;
		RECT	9.315 290.235 9.365 290.365 ;
		RECT	9.72 290.235 9.77 290.365 ;
		RECT	11.025 290.235 11.075 290.365 ;
		RECT	12.79 290.235 12.84 290.365 ;
		RECT	6.225 292.655 6.275 292.785 ;
		RECT	7.5 292.655 7.55 292.785 ;
		RECT	9.04 292.655 9.09 292.785 ;
		RECT	9.315 292.655 9.365 292.785 ;
		RECT	11.025 292.655 11.075 292.785 ;
		RECT	12.79 292.655 12.84 292.785 ;
		RECT	7.18 292.885 7.23 293.015 ;
		RECT	14.14 292.885 14.19 293.015 ;
		RECT	8.56 290.235 8.61 290.365 ;
		RECT	10.27 290.235 10.32 290.365 ;
		RECT	8.56 292.655 8.61 292.785 ;
		RECT	10.27 292.655 10.32 292.785 ;
		RECT	6.22 293.115 6.27 293.245 ;
		RECT	7.5 293.115 7.55 293.245 ;
		RECT	9.04 293.115 9.09 293.245 ;
		RECT	9.315 293.115 9.365 293.245 ;
		RECT	9.72 293.115 9.77 293.245 ;
		RECT	11.025 293.115 11.075 293.245 ;
		RECT	12.79 293.115 12.84 293.245 ;
		RECT	6.225 295.535 6.275 295.665 ;
		RECT	7.5 295.535 7.55 295.665 ;
		RECT	9.04 295.535 9.09 295.665 ;
		RECT	9.315 295.535 9.365 295.665 ;
		RECT	11.025 295.535 11.075 295.665 ;
		RECT	12.79 295.535 12.84 295.665 ;
		RECT	7.18 295.765 7.23 295.895 ;
		RECT	14.14 295.765 14.19 295.895 ;
		RECT	8.56 293.115 8.61 293.245 ;
		RECT	10.27 293.115 10.32 293.245 ;
		RECT	8.56 295.535 8.61 295.665 ;
		RECT	10.27 295.535 10.32 295.665 ;
		RECT	6.22 295.995 6.27 296.125 ;
		RECT	7.5 295.995 7.55 296.125 ;
		RECT	9.04 295.995 9.09 296.125 ;
		RECT	9.315 295.995 9.365 296.125 ;
		RECT	9.72 295.995 9.77 296.125 ;
		RECT	11.025 295.995 11.075 296.125 ;
		RECT	12.79 295.995 12.84 296.125 ;
		RECT	6.225 298.415 6.275 298.545 ;
		RECT	7.5 298.415 7.55 298.545 ;
		RECT	9.04 298.415 9.09 298.545 ;
		RECT	9.315 298.415 9.365 298.545 ;
		RECT	11.025 298.415 11.075 298.545 ;
		RECT	12.79 298.415 12.84 298.545 ;
		RECT	7.18 298.645 7.23 298.775 ;
		RECT	14.14 298.645 14.19 298.775 ;
		RECT	8.56 295.995 8.61 296.125 ;
		RECT	10.27 295.995 10.32 296.125 ;
		RECT	8.56 298.415 8.61 298.545 ;
		RECT	10.27 298.415 10.32 298.545 ;
		RECT	6.22 298.875 6.27 299.005 ;
		RECT	7.5 298.875 7.55 299.005 ;
		RECT	9.04 298.875 9.09 299.005 ;
		RECT	9.315 298.875 9.365 299.005 ;
		RECT	9.72 298.875 9.77 299.005 ;
		RECT	11.025 298.875 11.075 299.005 ;
		RECT	12.79 298.875 12.84 299.005 ;
		RECT	6.225 301.295 6.275 301.425 ;
		RECT	7.5 301.295 7.55 301.425 ;
		RECT	9.04 301.295 9.09 301.425 ;
		RECT	9.315 301.295 9.365 301.425 ;
		RECT	11.025 301.295 11.075 301.425 ;
		RECT	12.79 301.295 12.84 301.425 ;
		RECT	7.18 301.525 7.23 301.655 ;
		RECT	14.14 301.525 14.19 301.655 ;
		RECT	8.56 298.875 8.61 299.005 ;
		RECT	10.27 298.875 10.32 299.005 ;
		RECT	8.56 301.295 8.61 301.425 ;
		RECT	10.27 301.295 10.32 301.425 ;
		RECT	6.22 301.755 6.27 301.885 ;
		RECT	7.5 301.755 7.55 301.885 ;
		RECT	9.04 301.755 9.09 301.885 ;
		RECT	9.315 301.755 9.365 301.885 ;
		RECT	9.72 301.755 9.77 301.885 ;
		RECT	11.025 301.755 11.075 301.885 ;
		RECT	12.79 301.755 12.84 301.885 ;
		RECT	6.225 304.175 6.275 304.305 ;
		RECT	7.5 304.175 7.55 304.305 ;
		RECT	9.04 304.175 9.09 304.305 ;
		RECT	9.315 304.175 9.365 304.305 ;
		RECT	11.025 304.175 11.075 304.305 ;
		RECT	12.79 304.175 12.84 304.305 ;
		RECT	7.18 304.405 7.23 304.535 ;
		RECT	14.14 304.405 14.19 304.535 ;
		RECT	8.56 301.755 8.61 301.885 ;
		RECT	10.27 301.755 10.32 301.885 ;
		RECT	8.56 304.175 8.61 304.305 ;
		RECT	10.27 304.175 10.32 304.305 ;
		RECT	6.22 304.635 6.27 304.765 ;
		RECT	7.5 304.635 7.55 304.765 ;
		RECT	9.04 304.635 9.09 304.765 ;
		RECT	9.315 304.635 9.365 304.765 ;
		RECT	9.72 304.635 9.77 304.765 ;
		RECT	11.025 304.635 11.075 304.765 ;
		RECT	12.79 304.635 12.84 304.765 ;
		RECT	6.225 307.055 6.275 307.185 ;
		RECT	7.5 307.055 7.55 307.185 ;
		RECT	9.04 307.055 9.09 307.185 ;
		RECT	9.315 307.055 9.365 307.185 ;
		RECT	11.025 307.055 11.075 307.185 ;
		RECT	12.79 307.055 12.84 307.185 ;
		RECT	7.18 307.285 7.23 307.415 ;
		RECT	14.14 307.285 14.19 307.415 ;
		RECT	8.56 304.635 8.61 304.765 ;
		RECT	10.27 304.635 10.32 304.765 ;
		RECT	8.56 307.055 8.61 307.185 ;
		RECT	10.27 307.055 10.32 307.185 ;
		RECT	6.22 307.515 6.27 307.645 ;
		RECT	7.5 307.515 7.55 307.645 ;
		RECT	9.04 307.515 9.09 307.645 ;
		RECT	9.315 307.515 9.365 307.645 ;
		RECT	9.72 307.515 9.77 307.645 ;
		RECT	11.025 307.515 11.075 307.645 ;
		RECT	12.79 307.515 12.84 307.645 ;
		RECT	6.225 309.935 6.275 310.065 ;
		RECT	7.5 309.935 7.55 310.065 ;
		RECT	9.04 309.935 9.09 310.065 ;
		RECT	9.315 309.935 9.365 310.065 ;
		RECT	11.025 309.935 11.075 310.065 ;
		RECT	12.79 309.935 12.84 310.065 ;
		RECT	7.18 310.165 7.23 310.295 ;
		RECT	14.14 310.165 14.19 310.295 ;
		RECT	8.56 307.515 8.61 307.645 ;
		RECT	10.27 307.515 10.32 307.645 ;
		RECT	8.56 309.935 8.61 310.065 ;
		RECT	10.27 309.935 10.32 310.065 ;
		RECT	6.22 310.395 6.27 310.525 ;
		RECT	7.5 310.395 7.55 310.525 ;
		RECT	9.04 310.395 9.09 310.525 ;
		RECT	9.315 310.395 9.365 310.525 ;
		RECT	9.72 310.395 9.77 310.525 ;
		RECT	11.025 310.395 11.075 310.525 ;
		RECT	12.79 310.395 12.84 310.525 ;
		RECT	6.225 312.815 6.275 312.945 ;
		RECT	7.5 312.815 7.55 312.945 ;
		RECT	9.04 312.815 9.09 312.945 ;
		RECT	9.315 312.815 9.365 312.945 ;
		RECT	11.025 312.815 11.075 312.945 ;
		RECT	12.79 312.815 12.84 312.945 ;
		RECT	7.18 313.045 7.23 313.175 ;
		RECT	14.14 313.045 14.19 313.175 ;
		RECT	8.56 310.395 8.61 310.525 ;
		RECT	10.27 310.395 10.32 310.525 ;
		RECT	8.56 312.815 8.61 312.945 ;
		RECT	10.27 312.815 10.32 312.945 ;
		RECT	6.22 313.275 6.27 313.405 ;
		RECT	7.5 313.275 7.55 313.405 ;
		RECT	9.04 313.275 9.09 313.405 ;
		RECT	9.315 313.275 9.365 313.405 ;
		RECT	9.72 313.275 9.77 313.405 ;
		RECT	11.025 313.275 11.075 313.405 ;
		RECT	12.79 313.275 12.84 313.405 ;
		RECT	6.225 315.695 6.275 315.825 ;
		RECT	7.5 315.695 7.55 315.825 ;
		RECT	9.04 315.695 9.09 315.825 ;
		RECT	9.315 315.695 9.365 315.825 ;
		RECT	11.025 315.695 11.075 315.825 ;
		RECT	12.79 315.695 12.84 315.825 ;
		RECT	7.18 315.925 7.23 316.055 ;
		RECT	14.14 315.925 14.19 316.055 ;
		RECT	8.56 313.275 8.61 313.405 ;
		RECT	10.27 313.275 10.32 313.405 ;
		RECT	8.56 315.695 8.61 315.825 ;
		RECT	10.27 315.695 10.32 315.825 ;
		RECT	6.22 316.155 6.27 316.285 ;
		RECT	7.5 316.155 7.55 316.285 ;
		RECT	9.04 316.155 9.09 316.285 ;
		RECT	9.315 316.155 9.365 316.285 ;
		RECT	9.72 316.155 9.77 316.285 ;
		RECT	11.025 316.155 11.075 316.285 ;
		RECT	12.79 316.155 12.84 316.285 ;
		RECT	6.225 318.575 6.275 318.705 ;
		RECT	7.5 318.575 7.55 318.705 ;
		RECT	9.04 318.575 9.09 318.705 ;
		RECT	9.315 318.575 9.365 318.705 ;
		RECT	11.025 318.575 11.075 318.705 ;
		RECT	12.79 318.575 12.84 318.705 ;
		RECT	7.18 318.805 7.23 318.935 ;
		RECT	14.14 318.805 14.19 318.935 ;
		RECT	8.56 316.155 8.61 316.285 ;
		RECT	10.27 316.155 10.32 316.285 ;
		RECT	8.56 318.575 8.61 318.705 ;
		RECT	10.27 318.575 10.32 318.705 ;
		RECT	6.22 319.035 6.27 319.165 ;
		RECT	7.5 319.035 7.55 319.165 ;
		RECT	9.04 319.035 9.09 319.165 ;
		RECT	9.315 319.035 9.365 319.165 ;
		RECT	9.72 319.035 9.77 319.165 ;
		RECT	11.025 319.035 11.075 319.165 ;
		RECT	12.79 319.035 12.84 319.165 ;
		RECT	6.225 321.455 6.275 321.585 ;
		RECT	7.5 321.455 7.55 321.585 ;
		RECT	9.04 321.455 9.09 321.585 ;
		RECT	9.315 321.455 9.365 321.585 ;
		RECT	11.025 321.455 11.075 321.585 ;
		RECT	12.79 321.455 12.84 321.585 ;
		RECT	7.18 321.685 7.23 321.815 ;
		RECT	14.14 321.685 14.19 321.815 ;
		RECT	8.56 319.035 8.61 319.165 ;
		RECT	10.27 319.035 10.32 319.165 ;
		RECT	8.56 321.455 8.61 321.585 ;
		RECT	10.27 321.455 10.32 321.585 ;
		RECT	6.22 321.915 6.27 322.045 ;
		RECT	7.5 321.915 7.55 322.045 ;
		RECT	9.04 321.915 9.09 322.045 ;
		RECT	9.315 321.915 9.365 322.045 ;
		RECT	9.72 321.915 9.77 322.045 ;
		RECT	11.025 321.915 11.075 322.045 ;
		RECT	12.79 321.915 12.84 322.045 ;
		RECT	6.225 324.335 6.275 324.465 ;
		RECT	7.5 324.335 7.55 324.465 ;
		RECT	9.04 324.335 9.09 324.465 ;
		RECT	9.315 324.335 9.365 324.465 ;
		RECT	11.025 324.335 11.075 324.465 ;
		RECT	12.79 324.335 12.84 324.465 ;
		RECT	7.18 324.565 7.23 324.695 ;
		RECT	14.14 324.565 14.19 324.695 ;
		RECT	8.56 321.915 8.61 322.045 ;
		RECT	10.27 321.915 10.32 322.045 ;
		RECT	8.56 324.335 8.61 324.465 ;
		RECT	10.27 324.335 10.32 324.465 ;
		RECT	6.22 324.795 6.27 324.925 ;
		RECT	7.5 324.795 7.55 324.925 ;
		RECT	9.04 324.795 9.09 324.925 ;
		RECT	9.315 324.795 9.365 324.925 ;
		RECT	9.72 324.795 9.77 324.925 ;
		RECT	11.025 324.795 11.075 324.925 ;
		RECT	12.79 324.795 12.84 324.925 ;
		RECT	6.225 327.215 6.275 327.345 ;
		RECT	7.5 327.215 7.55 327.345 ;
		RECT	9.04 327.215 9.09 327.345 ;
		RECT	9.315 327.215 9.365 327.345 ;
		RECT	11.025 327.215 11.075 327.345 ;
		RECT	12.79 327.215 12.84 327.345 ;
		RECT	7.18 327.445 7.23 327.575 ;
		RECT	14.14 327.445 14.19 327.575 ;
		RECT	8.56 324.795 8.61 324.925 ;
		RECT	10.27 324.795 10.32 324.925 ;
		RECT	8.56 327.215 8.61 327.345 ;
		RECT	10.27 327.215 10.32 327.345 ;
		RECT	6.22 327.675 6.27 327.805 ;
		RECT	7.5 327.675 7.55 327.805 ;
		RECT	9.04 327.675 9.09 327.805 ;
		RECT	9.315 327.675 9.365 327.805 ;
		RECT	9.72 327.675 9.77 327.805 ;
		RECT	11.025 327.675 11.075 327.805 ;
		RECT	12.79 327.675 12.84 327.805 ;
		RECT	6.225 330.095 6.275 330.225 ;
		RECT	7.5 330.095 7.55 330.225 ;
		RECT	9.04 330.095 9.09 330.225 ;
		RECT	9.315 330.095 9.365 330.225 ;
		RECT	11.025 330.095 11.075 330.225 ;
		RECT	12.79 330.095 12.84 330.225 ;
		RECT	7.18 330.325 7.23 330.455 ;
		RECT	14.14 330.325 14.19 330.455 ;
		RECT	8.56 327.675 8.61 327.805 ;
		RECT	10.27 327.675 10.32 327.805 ;
		RECT	8.56 330.095 8.61 330.225 ;
		RECT	10.27 330.095 10.32 330.225 ;
		RECT	6.22 330.555 6.27 330.685 ;
		RECT	7.5 330.555 7.55 330.685 ;
		RECT	9.04 330.555 9.09 330.685 ;
		RECT	9.315 330.555 9.365 330.685 ;
		RECT	9.72 330.555 9.77 330.685 ;
		RECT	11.025 330.555 11.075 330.685 ;
		RECT	12.79 330.555 12.84 330.685 ;
		RECT	6.225 332.975 6.275 333.105 ;
		RECT	7.5 332.975 7.55 333.105 ;
		RECT	9.04 332.975 9.09 333.105 ;
		RECT	9.315 332.975 9.365 333.105 ;
		RECT	11.025 332.975 11.075 333.105 ;
		RECT	12.79 332.975 12.84 333.105 ;
		RECT	7.18 333.205 7.23 333.335 ;
		RECT	14.14 333.205 14.19 333.335 ;
		RECT	8.56 330.555 8.61 330.685 ;
		RECT	10.27 330.555 10.32 330.685 ;
		RECT	8.56 332.975 8.61 333.105 ;
		RECT	10.27 332.975 10.32 333.105 ;
		RECT	6.22 333.435 6.27 333.565 ;
		RECT	7.5 333.435 7.55 333.565 ;
		RECT	9.04 333.435 9.09 333.565 ;
		RECT	9.315 333.435 9.365 333.565 ;
		RECT	9.72 333.435 9.77 333.565 ;
		RECT	11.025 333.435 11.075 333.565 ;
		RECT	12.79 333.435 12.84 333.565 ;
		RECT	6.225 335.855 6.275 335.985 ;
		RECT	7.5 335.855 7.55 335.985 ;
		RECT	9.04 335.855 9.09 335.985 ;
		RECT	9.315 335.855 9.365 335.985 ;
		RECT	11.025 335.855 11.075 335.985 ;
		RECT	12.79 335.855 12.84 335.985 ;
		RECT	7.18 336.085 7.23 336.215 ;
		RECT	14.14 336.085 14.19 336.215 ;
		RECT	8.56 333.435 8.61 333.565 ;
		RECT	10.27 333.435 10.32 333.565 ;
		RECT	8.56 335.855 8.61 335.985 ;
		RECT	10.27 335.855 10.32 335.985 ;
		RECT	6.22 336.315 6.27 336.445 ;
		RECT	7.5 336.315 7.55 336.445 ;
		RECT	9.04 336.315 9.09 336.445 ;
		RECT	9.315 336.315 9.365 336.445 ;
		RECT	9.72 336.315 9.77 336.445 ;
		RECT	11.025 336.315 11.075 336.445 ;
		RECT	12.79 336.315 12.84 336.445 ;
		RECT	6.225 338.735 6.275 338.865 ;
		RECT	7.5 338.735 7.55 338.865 ;
		RECT	9.04 338.735 9.09 338.865 ;
		RECT	9.315 338.735 9.365 338.865 ;
		RECT	11.025 338.735 11.075 338.865 ;
		RECT	12.79 338.735 12.84 338.865 ;
		RECT	7.18 338.965 7.23 339.095 ;
		RECT	14.14 338.965 14.19 339.095 ;
		RECT	8.56 336.315 8.61 336.445 ;
		RECT	10.27 336.315 10.32 336.445 ;
		RECT	8.56 338.735 8.61 338.865 ;
		RECT	10.27 338.735 10.32 338.865 ;
		RECT	6.22 339.195 6.27 339.325 ;
		RECT	7.5 339.195 7.55 339.325 ;
		RECT	9.04 339.195 9.09 339.325 ;
		RECT	9.315 339.195 9.365 339.325 ;
		RECT	9.72 339.195 9.77 339.325 ;
		RECT	11.025 339.195 11.075 339.325 ;
		RECT	12.79 339.195 12.84 339.325 ;
		RECT	6.225 341.615 6.275 341.745 ;
		RECT	7.5 341.615 7.55 341.745 ;
		RECT	9.04 341.615 9.09 341.745 ;
		RECT	9.315 341.615 9.365 341.745 ;
		RECT	11.025 341.615 11.075 341.745 ;
		RECT	12.79 341.615 12.84 341.745 ;
		RECT	7.18 341.845 7.23 341.975 ;
		RECT	14.14 341.845 14.19 341.975 ;
		RECT	8.56 339.195 8.61 339.325 ;
		RECT	10.27 339.195 10.32 339.325 ;
		RECT	8.56 341.615 8.61 341.745 ;
		RECT	10.27 341.615 10.32 341.745 ;
		RECT	6.22 342.075 6.27 342.205 ;
		RECT	7.5 342.075 7.55 342.205 ;
		RECT	9.04 342.075 9.09 342.205 ;
		RECT	9.315 342.075 9.365 342.205 ;
		RECT	9.72 342.075 9.77 342.205 ;
		RECT	11.025 342.075 11.075 342.205 ;
		RECT	12.79 342.075 12.84 342.205 ;
		RECT	6.225 344.495 6.275 344.625 ;
		RECT	7.5 344.495 7.55 344.625 ;
		RECT	9.04 344.495 9.09 344.625 ;
		RECT	9.315 344.495 9.365 344.625 ;
		RECT	11.025 344.495 11.075 344.625 ;
		RECT	12.79 344.495 12.84 344.625 ;
		RECT	7.18 344.725 7.23 344.855 ;
		RECT	14.14 344.725 14.19 344.855 ;
		RECT	8.56 342.075 8.61 342.205 ;
		RECT	10.27 342.075 10.32 342.205 ;
		RECT	8.56 344.495 8.61 344.625 ;
		RECT	10.27 344.495 10.32 344.625 ;
		RECT	6.22 344.955 6.27 345.085 ;
		RECT	7.5 344.955 7.55 345.085 ;
		RECT	9.04 344.955 9.09 345.085 ;
		RECT	9.315 344.955 9.365 345.085 ;
		RECT	9.72 344.955 9.77 345.085 ;
		RECT	11.025 344.955 11.075 345.085 ;
		RECT	12.79 344.955 12.84 345.085 ;
		RECT	6.225 347.375 6.275 347.505 ;
		RECT	7.5 347.375 7.55 347.505 ;
		RECT	9.04 347.375 9.09 347.505 ;
		RECT	9.315 347.375 9.365 347.505 ;
		RECT	11.025 347.375 11.075 347.505 ;
		RECT	12.79 347.375 12.84 347.505 ;
		RECT	7.18 347.605 7.23 347.735 ;
		RECT	14.14 347.605 14.19 347.735 ;
		RECT	8.56 344.955 8.61 345.085 ;
		RECT	10.27 344.955 10.32 345.085 ;
		RECT	8.56 347.375 8.61 347.505 ;
		RECT	10.27 347.375 10.32 347.505 ;
		RECT	6.22 347.835 6.27 347.965 ;
		RECT	7.5 347.835 7.55 347.965 ;
		RECT	9.04 347.835 9.09 347.965 ;
		RECT	9.315 347.835 9.365 347.965 ;
		RECT	9.72 347.835 9.77 347.965 ;
		RECT	11.025 347.835 11.075 347.965 ;
		RECT	12.79 347.835 12.84 347.965 ;
		RECT	6.225 350.255 6.275 350.385 ;
		RECT	7.5 350.255 7.55 350.385 ;
		RECT	9.04 350.255 9.09 350.385 ;
		RECT	9.315 350.255 9.365 350.385 ;
		RECT	11.025 350.255 11.075 350.385 ;
		RECT	12.79 350.255 12.84 350.385 ;
		RECT	7.18 350.485 7.23 350.615 ;
		RECT	14.14 350.485 14.19 350.615 ;
		RECT	8.56 347.835 8.61 347.965 ;
		RECT	10.27 347.835 10.32 347.965 ;
		RECT	8.56 350.255 8.61 350.385 ;
		RECT	10.27 350.255 10.32 350.385 ;
		RECT	6.22 350.715 6.27 350.845 ;
		RECT	7.5 350.715 7.55 350.845 ;
		RECT	9.04 350.715 9.09 350.845 ;
		RECT	9.315 350.715 9.365 350.845 ;
		RECT	9.72 350.715 9.77 350.845 ;
		RECT	11.025 350.715 11.075 350.845 ;
		RECT	12.79 350.715 12.84 350.845 ;
		RECT	6.225 353.135 6.275 353.265 ;
		RECT	7.5 353.135 7.55 353.265 ;
		RECT	9.04 353.135 9.09 353.265 ;
		RECT	9.315 353.135 9.365 353.265 ;
		RECT	11.025 353.135 11.075 353.265 ;
		RECT	12.79 353.135 12.84 353.265 ;
		RECT	7.18 353.365 7.23 353.495 ;
		RECT	14.14 353.365 14.19 353.495 ;
		RECT	8.56 350.715 8.61 350.845 ;
		RECT	10.27 350.715 10.32 350.845 ;
		RECT	8.56 353.135 8.61 353.265 ;
		RECT	10.27 353.135 10.32 353.265 ;
		RECT	6.22 353.595 6.27 353.725 ;
		RECT	7.5 353.595 7.55 353.725 ;
		RECT	9.04 353.595 9.09 353.725 ;
		RECT	9.315 353.595 9.365 353.725 ;
		RECT	9.72 353.595 9.77 353.725 ;
		RECT	11.025 353.595 11.075 353.725 ;
		RECT	12.79 353.595 12.84 353.725 ;
		RECT	6.225 356.015 6.275 356.145 ;
		RECT	7.5 356.015 7.55 356.145 ;
		RECT	9.04 356.015 9.09 356.145 ;
		RECT	9.315 356.015 9.365 356.145 ;
		RECT	11.025 356.015 11.075 356.145 ;
		RECT	12.79 356.015 12.84 356.145 ;
		RECT	7.18 356.245 7.23 356.375 ;
		RECT	14.14 356.245 14.19 356.375 ;
		RECT	8.56 353.595 8.61 353.725 ;
		RECT	10.27 353.595 10.32 353.725 ;
		RECT	8.56 356.015 8.61 356.145 ;
		RECT	10.27 356.015 10.32 356.145 ;
		RECT	6.22 356.475 6.27 356.605 ;
		RECT	7.5 356.475 7.55 356.605 ;
		RECT	9.04 356.475 9.09 356.605 ;
		RECT	9.315 356.475 9.365 356.605 ;
		RECT	9.72 356.475 9.77 356.605 ;
		RECT	11.025 356.475 11.075 356.605 ;
		RECT	12.79 356.475 12.84 356.605 ;
		RECT	6.225 358.895 6.275 359.025 ;
		RECT	7.5 358.895 7.55 359.025 ;
		RECT	9.04 358.895 9.09 359.025 ;
		RECT	9.315 358.895 9.365 359.025 ;
		RECT	11.025 358.895 11.075 359.025 ;
		RECT	12.79 358.895 12.84 359.025 ;
		RECT	7.18 359.125 7.23 359.255 ;
		RECT	14.14 359.125 14.19 359.255 ;
		RECT	8.56 356.475 8.61 356.605 ;
		RECT	10.27 356.475 10.32 356.605 ;
		RECT	8.56 358.895 8.61 359.025 ;
		RECT	10.27 358.895 10.32 359.025 ;
		RECT	6.22 359.355 6.27 359.485 ;
		RECT	7.5 359.355 7.55 359.485 ;
		RECT	9.04 359.355 9.09 359.485 ;
		RECT	9.315 359.355 9.365 359.485 ;
		RECT	9.72 359.355 9.77 359.485 ;
		RECT	11.025 359.355 11.075 359.485 ;
		RECT	12.79 359.355 12.84 359.485 ;
		RECT	6.225 361.775 6.275 361.905 ;
		RECT	7.5 361.775 7.55 361.905 ;
		RECT	9.04 361.775 9.09 361.905 ;
		RECT	9.315 361.775 9.365 361.905 ;
		RECT	11.025 361.775 11.075 361.905 ;
		RECT	12.79 361.775 12.84 361.905 ;
		RECT	7.18 362.005 7.23 362.135 ;
		RECT	14.14 362.005 14.19 362.135 ;
		RECT	8.56 359.355 8.61 359.485 ;
		RECT	10.27 359.355 10.32 359.485 ;
		RECT	8.56 361.775 8.61 361.905 ;
		RECT	10.27 361.775 10.32 361.905 ;
		RECT	6.22 362.235 6.27 362.365 ;
		RECT	7.5 362.235 7.55 362.365 ;
		RECT	9.04 362.235 9.09 362.365 ;
		RECT	9.315 362.235 9.365 362.365 ;
		RECT	9.72 362.235 9.77 362.365 ;
		RECT	11.025 362.235 11.075 362.365 ;
		RECT	12.79 362.235 12.84 362.365 ;
		RECT	6.225 364.655 6.275 364.785 ;
		RECT	7.5 364.655 7.55 364.785 ;
		RECT	9.04 364.655 9.09 364.785 ;
		RECT	9.315 364.655 9.365 364.785 ;
		RECT	11.025 364.655 11.075 364.785 ;
		RECT	12.79 364.655 12.84 364.785 ;
		RECT	7.18 364.885 7.23 365.015 ;
		RECT	14.14 364.885 14.19 365.015 ;
		RECT	8.56 362.235 8.61 362.365 ;
		RECT	10.27 362.235 10.32 362.365 ;
		RECT	8.56 364.655 8.61 364.785 ;
		RECT	10.27 364.655 10.32 364.785 ;
		RECT	6.22 365.115 6.27 365.245 ;
		RECT	7.5 365.115 7.55 365.245 ;
		RECT	9.04 365.115 9.09 365.245 ;
		RECT	9.315 365.115 9.365 365.245 ;
		RECT	9.72 365.115 9.77 365.245 ;
		RECT	11.025 365.115 11.075 365.245 ;
		RECT	12.79 365.115 12.84 365.245 ;
		RECT	6.225 367.535 6.275 367.665 ;
		RECT	7.5 367.535 7.55 367.665 ;
		RECT	9.04 367.535 9.09 367.665 ;
		RECT	9.315 367.535 9.365 367.665 ;
		RECT	11.025 367.535 11.075 367.665 ;
		RECT	12.79 367.535 12.84 367.665 ;
		RECT	7.18 367.765 7.23 367.895 ;
		RECT	14.14 367.765 14.19 367.895 ;
		RECT	8.56 365.115 8.61 365.245 ;
		RECT	10.27 365.115 10.32 365.245 ;
		RECT	8.56 367.535 8.61 367.665 ;
		RECT	10.27 367.535 10.32 367.665 ;
		RECT	6.22 367.995 6.27 368.125 ;
		RECT	7.5 367.995 7.55 368.125 ;
		RECT	9.04 367.995 9.09 368.125 ;
		RECT	9.315 367.995 9.365 368.125 ;
		RECT	9.72 367.995 9.77 368.125 ;
		RECT	11.025 367.995 11.075 368.125 ;
		RECT	12.79 367.995 12.84 368.125 ;
		RECT	6.225 370.415 6.275 370.545 ;
		RECT	7.5 370.415 7.55 370.545 ;
		RECT	9.04 370.415 9.09 370.545 ;
		RECT	9.315 370.415 9.365 370.545 ;
		RECT	11.025 370.415 11.075 370.545 ;
		RECT	12.79 370.415 12.84 370.545 ;
		RECT	7.18 370.645 7.23 370.775 ;
		RECT	14.14 370.645 14.19 370.775 ;
		RECT	8.56 367.995 8.61 368.125 ;
		RECT	10.27 367.995 10.32 368.125 ;
		RECT	8.56 370.415 8.61 370.545 ;
		RECT	10.27 370.415 10.32 370.545 ;
		RECT	6.22 370.875 6.27 371.005 ;
		RECT	7.5 370.875 7.55 371.005 ;
		RECT	9.04 370.875 9.09 371.005 ;
		RECT	9.315 370.875 9.365 371.005 ;
		RECT	9.72 370.875 9.77 371.005 ;
		RECT	11.025 370.875 11.075 371.005 ;
		RECT	12.79 370.875 12.84 371.005 ;
		RECT	6.225 373.295 6.275 373.425 ;
		RECT	7.5 373.295 7.55 373.425 ;
		RECT	9.04 373.295 9.09 373.425 ;
		RECT	9.315 373.295 9.365 373.425 ;
		RECT	11.025 373.295 11.075 373.425 ;
		RECT	12.79 373.295 12.84 373.425 ;
		RECT	7.18 373.525 7.23 373.655 ;
		RECT	14.14 373.525 14.19 373.655 ;
		RECT	8.56 370.875 8.61 371.005 ;
		RECT	10.27 370.875 10.32 371.005 ;
		RECT	8.56 373.295 8.61 373.425 ;
		RECT	10.27 373.295 10.32 373.425 ;
		RECT	6.22 373.755 6.27 373.885 ;
		RECT	7.5 373.755 7.55 373.885 ;
		RECT	9.04 373.755 9.09 373.885 ;
		RECT	9.315 373.755 9.365 373.885 ;
		RECT	9.72 373.755 9.77 373.885 ;
		RECT	11.025 373.755 11.075 373.885 ;
		RECT	12.79 373.755 12.84 373.885 ;
		RECT	6.225 376.175 6.275 376.305 ;
		RECT	7.5 376.175 7.55 376.305 ;
		RECT	9.04 376.175 9.09 376.305 ;
		RECT	9.315 376.175 9.365 376.305 ;
		RECT	11.025 376.175 11.075 376.305 ;
		RECT	12.79 376.175 12.84 376.305 ;
		RECT	7.18 376.405 7.23 376.535 ;
		RECT	14.14 376.405 14.19 376.535 ;
		RECT	8.56 373.755 8.61 373.885 ;
		RECT	10.27 373.755 10.32 373.885 ;
		RECT	8.56 376.175 8.61 376.305 ;
		RECT	10.27 376.175 10.32 376.305 ;
		RECT	6.22 376.635 6.27 376.765 ;
		RECT	7.5 376.635 7.55 376.765 ;
		RECT	9.04 376.635 9.09 376.765 ;
		RECT	9.315 376.635 9.365 376.765 ;
		RECT	9.72 376.635 9.77 376.765 ;
		RECT	11.025 376.635 11.075 376.765 ;
		RECT	12.79 376.635 12.84 376.765 ;
		RECT	6.225 379.055 6.275 379.185 ;
		RECT	7.5 379.055 7.55 379.185 ;
		RECT	9.04 379.055 9.09 379.185 ;
		RECT	9.315 379.055 9.365 379.185 ;
		RECT	11.025 379.055 11.075 379.185 ;
		RECT	12.79 379.055 12.84 379.185 ;
		RECT	7.18 379.285 7.23 379.415 ;
		RECT	14.14 379.285 14.19 379.415 ;
		RECT	8.56 376.635 8.61 376.765 ;
		RECT	10.27 376.635 10.32 376.765 ;
		RECT	8.56 379.055 8.61 379.185 ;
		RECT	10.27 379.055 10.32 379.185 ;
		RECT	6.22 379.515 6.27 379.645 ;
		RECT	7.5 379.515 7.55 379.645 ;
		RECT	9.04 379.515 9.09 379.645 ;
		RECT	9.315 379.515 9.365 379.645 ;
		RECT	9.72 379.515 9.77 379.645 ;
		RECT	11.025 379.515 11.075 379.645 ;
		RECT	12.79 379.515 12.84 379.645 ;
		RECT	6.225 381.935 6.275 382.065 ;
		RECT	7.5 381.935 7.55 382.065 ;
		RECT	9.04 381.935 9.09 382.065 ;
		RECT	9.315 381.935 9.365 382.065 ;
		RECT	11.025 381.935 11.075 382.065 ;
		RECT	12.79 381.935 12.84 382.065 ;
		RECT	7.18 382.165 7.23 382.295 ;
		RECT	14.14 382.165 14.19 382.295 ;
		RECT	8.56 379.515 8.61 379.645 ;
		RECT	10.27 379.515 10.32 379.645 ;
		RECT	8.56 381.935 8.61 382.065 ;
		RECT	10.27 381.935 10.32 382.065 ;
		RECT	6.22 382.395 6.27 382.525 ;
		RECT	7.5 382.395 7.55 382.525 ;
		RECT	9.04 382.395 9.09 382.525 ;
		RECT	9.315 382.395 9.365 382.525 ;
		RECT	9.72 382.395 9.77 382.525 ;
		RECT	11.025 382.395 11.075 382.525 ;
		RECT	12.79 382.395 12.84 382.525 ;
		RECT	6.225 384.815 6.275 384.945 ;
		RECT	7.5 384.815 7.55 384.945 ;
		RECT	9.04 384.815 9.09 384.945 ;
		RECT	9.315 384.815 9.365 384.945 ;
		RECT	11.025 384.815 11.075 384.945 ;
		RECT	12.79 384.815 12.84 384.945 ;
		RECT	7.18 385.045 7.23 385.175 ;
		RECT	14.14 385.045 14.19 385.175 ;
		RECT	8.56 382.395 8.61 382.525 ;
		RECT	10.27 382.395 10.32 382.525 ;
		RECT	8.56 384.815 8.61 384.945 ;
		RECT	10.27 384.815 10.32 384.945 ;
		RECT	6.22 385.275 6.27 385.405 ;
		RECT	7.5 385.275 7.55 385.405 ;
		RECT	9.04 385.275 9.09 385.405 ;
		RECT	9.315 385.275 9.365 385.405 ;
		RECT	9.72 385.275 9.77 385.405 ;
		RECT	11.025 385.275 11.075 385.405 ;
		RECT	12.79 385.275 12.84 385.405 ;
		RECT	6.225 387.695 6.275 387.825 ;
		RECT	7.5 387.695 7.55 387.825 ;
		RECT	9.04 387.695 9.09 387.825 ;
		RECT	9.315 387.695 9.365 387.825 ;
		RECT	11.025 387.695 11.075 387.825 ;
		RECT	12.79 387.695 12.84 387.825 ;
		RECT	7.18 387.925 7.23 388.055 ;
		RECT	14.14 387.925 14.19 388.055 ;
		RECT	8.56 385.275 8.61 385.405 ;
		RECT	10.27 385.275 10.32 385.405 ;
		RECT	8.56 387.695 8.61 387.825 ;
		RECT	10.27 387.695 10.32 387.825 ;
		RECT	6.22 388.155 6.27 388.285 ;
		RECT	7.5 388.155 7.55 388.285 ;
		RECT	9.04 388.155 9.09 388.285 ;
		RECT	9.315 388.155 9.365 388.285 ;
		RECT	9.72 388.155 9.77 388.285 ;
		RECT	11.025 388.155 11.075 388.285 ;
		RECT	12.79 388.155 12.84 388.285 ;
		RECT	6.225 390.575 6.275 390.705 ;
		RECT	7.5 390.575 7.55 390.705 ;
		RECT	9.04 390.575 9.09 390.705 ;
		RECT	9.315 390.575 9.365 390.705 ;
		RECT	11.025 390.575 11.075 390.705 ;
		RECT	12.79 390.575 12.84 390.705 ;
		RECT	7.18 390.805 7.23 390.935 ;
		RECT	14.14 390.805 14.19 390.935 ;
		RECT	8.56 388.155 8.61 388.285 ;
		RECT	10.27 388.155 10.32 388.285 ;
		RECT	8.56 390.575 8.61 390.705 ;
		RECT	10.27 390.575 10.32 390.705 ;
		RECT	6.22 391.035 6.27 391.165 ;
		RECT	7.5 391.035 7.55 391.165 ;
		RECT	9.04 391.035 9.09 391.165 ;
		RECT	9.315 391.035 9.365 391.165 ;
		RECT	9.72 391.035 9.77 391.165 ;
		RECT	11.025 391.035 11.075 391.165 ;
		RECT	12.79 391.035 12.84 391.165 ;
		RECT	6.225 393.455 6.275 393.585 ;
		RECT	7.5 393.455 7.55 393.585 ;
		RECT	9.04 393.455 9.09 393.585 ;
		RECT	9.315 393.455 9.365 393.585 ;
		RECT	11.025 393.455 11.075 393.585 ;
		RECT	12.79 393.455 12.84 393.585 ;
		RECT	7.18 393.685 7.23 393.815 ;
		RECT	14.14 393.685 14.19 393.815 ;
		RECT	8.56 391.035 8.61 391.165 ;
		RECT	10.27 391.035 10.32 391.165 ;
		RECT	8.56 393.455 8.61 393.585 ;
		RECT	10.27 393.455 10.32 393.585 ;
		RECT	6.22 393.915 6.27 394.045 ;
		RECT	7.5 393.915 7.55 394.045 ;
		RECT	9.04 393.915 9.09 394.045 ;
		RECT	9.315 393.915 9.365 394.045 ;
		RECT	9.72 393.915 9.77 394.045 ;
		RECT	11.025 393.915 11.075 394.045 ;
		RECT	12.79 393.915 12.84 394.045 ;
		RECT	6.225 396.335 6.275 396.465 ;
		RECT	7.5 396.335 7.55 396.465 ;
		RECT	9.04 396.335 9.09 396.465 ;
		RECT	9.315 396.335 9.365 396.465 ;
		RECT	11.025 396.335 11.075 396.465 ;
		RECT	12.79 396.335 12.84 396.465 ;
		RECT	7.18 396.565 7.23 396.695 ;
		RECT	14.14 396.565 14.19 396.695 ;
		RECT	8.56 393.915 8.61 394.045 ;
		RECT	10.27 393.915 10.32 394.045 ;
		RECT	8.56 396.335 8.61 396.465 ;
		RECT	10.27 396.335 10.32 396.465 ;
		RECT	6.22 396.795 6.27 396.925 ;
		RECT	7.5 396.795 7.55 396.925 ;
		RECT	9.04 396.795 9.09 396.925 ;
		RECT	9.315 396.795 9.365 396.925 ;
		RECT	9.72 396.795 9.77 396.925 ;
		RECT	11.025 396.795 11.075 396.925 ;
		RECT	12.79 396.795 12.84 396.925 ;
		RECT	6.225 399.215 6.275 399.345 ;
		RECT	7.5 399.215 7.55 399.345 ;
		RECT	9.04 399.215 9.09 399.345 ;
		RECT	9.315 399.215 9.365 399.345 ;
		RECT	11.025 399.215 11.075 399.345 ;
		RECT	12.79 399.215 12.84 399.345 ;
		RECT	7.18 399.445 7.23 399.575 ;
		RECT	14.14 399.445 14.19 399.575 ;
		RECT	8.56 396.795 8.61 396.925 ;
		RECT	10.27 396.795 10.32 396.925 ;
		RECT	8.56 399.215 8.61 399.345 ;
		RECT	10.27 399.215 10.32 399.345 ;
		RECT	6.22 399.675 6.27 399.805 ;
		RECT	7.5 399.675 7.55 399.805 ;
		RECT	9.04 399.675 9.09 399.805 ;
		RECT	9.315 399.675 9.365 399.805 ;
		RECT	9.72 399.675 9.77 399.805 ;
		RECT	11.025 399.675 11.075 399.805 ;
		RECT	12.79 399.675 12.84 399.805 ;
		RECT	6.225 402.095 6.275 402.225 ;
		RECT	7.5 402.095 7.55 402.225 ;
		RECT	9.04 402.095 9.09 402.225 ;
		RECT	9.315 402.095 9.365 402.225 ;
		RECT	11.025 402.095 11.075 402.225 ;
		RECT	12.79 402.095 12.84 402.225 ;
		RECT	7.18 402.325 7.23 402.455 ;
		RECT	14.14 402.325 14.19 402.455 ;
		RECT	8.56 399.675 8.61 399.805 ;
		RECT	10.27 399.675 10.32 399.805 ;
		RECT	8.56 402.095 8.61 402.225 ;
		RECT	10.27 402.095 10.32 402.225 ;
		RECT	6.22 402.555 6.27 402.685 ;
		RECT	7.5 402.555 7.55 402.685 ;
		RECT	9.04 402.555 9.09 402.685 ;
		RECT	9.315 402.555 9.365 402.685 ;
		RECT	9.72 402.555 9.77 402.685 ;
		RECT	11.025 402.555 11.075 402.685 ;
		RECT	12.79 402.555 12.84 402.685 ;
		RECT	6.225 404.975 6.275 405.105 ;
		RECT	7.5 404.975 7.55 405.105 ;
		RECT	9.04 404.975 9.09 405.105 ;
		RECT	9.315 404.975 9.365 405.105 ;
		RECT	11.025 404.975 11.075 405.105 ;
		RECT	12.79 404.975 12.84 405.105 ;
		RECT	7.18 405.205 7.23 405.335 ;
		RECT	14.14 405.205 14.19 405.335 ;
		RECT	8.56 402.555 8.61 402.685 ;
		RECT	10.27 402.555 10.32 402.685 ;
		RECT	8.56 404.975 8.61 405.105 ;
		RECT	10.27 404.975 10.32 405.105 ;
		RECT	6.22 405.435 6.27 405.565 ;
		RECT	7.5 405.435 7.55 405.565 ;
		RECT	9.04 405.435 9.09 405.565 ;
		RECT	9.315 405.435 9.365 405.565 ;
		RECT	9.72 405.435 9.77 405.565 ;
		RECT	11.025 405.435 11.075 405.565 ;
		RECT	12.79 405.435 12.84 405.565 ;
		RECT	6.225 407.855 6.275 407.985 ;
		RECT	7.5 407.855 7.55 407.985 ;
		RECT	9.04 407.855 9.09 407.985 ;
		RECT	9.315 407.855 9.365 407.985 ;
		RECT	11.025 407.855 11.075 407.985 ;
		RECT	12.79 407.855 12.84 407.985 ;
		RECT	7.18 408.085 7.23 408.215 ;
		RECT	14.14 408.085 14.19 408.215 ;
		RECT	8.56 405.435 8.61 405.565 ;
		RECT	10.27 405.435 10.32 405.565 ;
		RECT	8.56 407.855 8.61 407.985 ;
		RECT	10.27 407.855 10.32 407.985 ;
		RECT	6.22 408.315 6.27 408.445 ;
		RECT	7.5 408.315 7.55 408.445 ;
		RECT	9.04 408.315 9.09 408.445 ;
		RECT	9.315 408.315 9.365 408.445 ;
		RECT	9.72 408.315 9.77 408.445 ;
		RECT	11.025 408.315 11.075 408.445 ;
		RECT	12.79 408.315 12.84 408.445 ;
		RECT	6.225 410.735 6.275 410.865 ;
		RECT	7.5 410.735 7.55 410.865 ;
		RECT	9.04 410.735 9.09 410.865 ;
		RECT	9.315 410.735 9.365 410.865 ;
		RECT	11.025 410.735 11.075 410.865 ;
		RECT	12.79 410.735 12.84 410.865 ;
		RECT	7.18 410.965 7.23 411.095 ;
		RECT	14.14 410.965 14.19 411.095 ;
		RECT	8.56 408.315 8.61 408.445 ;
		RECT	10.27 408.315 10.32 408.445 ;
		RECT	8.56 410.735 8.61 410.865 ;
		RECT	10.27 410.735 10.32 410.865 ;
		RECT	6.22 411.195 6.27 411.325 ;
		RECT	7.5 411.195 7.55 411.325 ;
		RECT	9.04 411.195 9.09 411.325 ;
		RECT	9.315 411.195 9.365 411.325 ;
		RECT	9.72 411.195 9.77 411.325 ;
		RECT	11.025 411.195 11.075 411.325 ;
		RECT	12.79 411.195 12.84 411.325 ;
		RECT	6.225 413.615 6.275 413.745 ;
		RECT	7.5 413.615 7.55 413.745 ;
		RECT	9.04 413.615 9.09 413.745 ;
		RECT	9.315 413.615 9.365 413.745 ;
		RECT	11.025 413.615 11.075 413.745 ;
		RECT	12.79 413.615 12.84 413.745 ;
		RECT	7.18 413.845 7.23 413.975 ;
		RECT	14.14 413.845 14.19 413.975 ;
		RECT	8.56 411.195 8.61 411.325 ;
		RECT	10.27 411.195 10.32 411.325 ;
		RECT	8.56 413.615 8.61 413.745 ;
		RECT	10.27 413.615 10.32 413.745 ;
		RECT	14.33 232.635 14.38 232.765 ;
		RECT	6.22 233.095 6.27 233.225 ;
		RECT	7.5 233.095 7.55 233.225 ;
		RECT	9.04 233.095 9.09 233.225 ;
		RECT	9.315 233.095 9.365 233.225 ;
		RECT	9.72 233.095 9.77 233.225 ;
		RECT	11.025 233.095 11.075 233.225 ;
		RECT	12.79 233.095 12.84 233.225 ;
		RECT	14.33 235.055 14.38 235.185 ;
		RECT	5.675 235.285 5.725 235.415 ;
		RECT	6.065 235.285 6.115 235.415 ;
		RECT	6.725 235.285 6.775 235.415 ;
		RECT	8.42 235.285 8.47 235.415 ;
		RECT	8.77 235.285 8.82 235.415 ;
		RECT	11.555 235.285 11.605 235.415 ;
		RECT	11.815 235.285 11.865 235.415 ;
		RECT	12.52 235.285 12.57 235.415 ;
		RECT	13.98 235.285 14.03 235.415 ;
		RECT	14.33 258.555 14.38 258.685 ;
		RECT	6.22 259.015 6.27 259.145 ;
		RECT	7.5 259.015 7.55 259.145 ;
		RECT	9.04 259.015 9.09 259.145 ;
		RECT	9.315 259.015 9.365 259.145 ;
		RECT	9.72 259.015 9.77 259.145 ;
		RECT	11.025 259.015 11.075 259.145 ;
		RECT	12.79 259.015 12.84 259.145 ;
		RECT	14.33 260.975 14.38 261.105 ;
		RECT	5.675 261.205 5.725 261.335 ;
		RECT	6.065 261.205 6.115 261.335 ;
		RECT	6.725 261.205 6.775 261.335 ;
		RECT	8.42 261.205 8.47 261.335 ;
		RECT	8.77 261.205 8.82 261.335 ;
		RECT	11.555 261.205 11.605 261.335 ;
		RECT	11.815 261.205 11.865 261.335 ;
		RECT	12.52 261.205 12.57 261.335 ;
		RECT	13.98 261.205 14.03 261.335 ;
		RECT	14.33 261.435 14.38 261.565 ;
		RECT	6.22 261.895 6.27 262.025 ;
		RECT	7.5 261.895 7.55 262.025 ;
		RECT	9.04 261.895 9.09 262.025 ;
		RECT	9.315 261.895 9.365 262.025 ;
		RECT	9.72 261.895 9.77 262.025 ;
		RECT	11.025 261.895 11.075 262.025 ;
		RECT	12.79 261.895 12.84 262.025 ;
		RECT	14.33 263.855 14.38 263.985 ;
		RECT	5.675 264.085 5.725 264.215 ;
		RECT	6.065 264.085 6.115 264.215 ;
		RECT	6.725 264.085 6.775 264.215 ;
		RECT	8.42 264.085 8.47 264.215 ;
		RECT	8.77 264.085 8.82 264.215 ;
		RECT	11.555 264.085 11.605 264.215 ;
		RECT	11.815 264.085 11.865 264.215 ;
		RECT	12.52 264.085 12.57 264.215 ;
		RECT	13.98 264.085 14.03 264.215 ;
		RECT	14.33 264.315 14.38 264.445 ;
		RECT	6.22 264.775 6.27 264.905 ;
		RECT	7.5 264.775 7.55 264.905 ;
		RECT	9.04 264.775 9.09 264.905 ;
		RECT	9.315 264.775 9.365 264.905 ;
		RECT	9.72 264.775 9.77 264.905 ;
		RECT	11.025 264.775 11.075 264.905 ;
		RECT	12.79 264.775 12.84 264.905 ;
		RECT	14.33 266.735 14.38 266.865 ;
		RECT	5.675 266.965 5.725 267.095 ;
		RECT	6.065 266.965 6.115 267.095 ;
		RECT	6.725 266.965 6.775 267.095 ;
		RECT	8.42 266.965 8.47 267.095 ;
		RECT	8.77 266.965 8.82 267.095 ;
		RECT	11.555 266.965 11.605 267.095 ;
		RECT	11.815 266.965 11.865 267.095 ;
		RECT	12.52 266.965 12.57 267.095 ;
		RECT	13.98 266.965 14.03 267.095 ;
		RECT	14.33 267.195 14.38 267.325 ;
		RECT	6.22 267.655 6.27 267.785 ;
		RECT	7.5 267.655 7.55 267.785 ;
		RECT	9.04 267.655 9.09 267.785 ;
		RECT	9.315 267.655 9.365 267.785 ;
		RECT	9.72 267.655 9.77 267.785 ;
		RECT	11.025 267.655 11.075 267.785 ;
		RECT	12.79 267.655 12.84 267.785 ;
		RECT	14.33 269.615 14.38 269.745 ;
		RECT	5.675 269.845 5.725 269.975 ;
		RECT	6.065 269.845 6.115 269.975 ;
		RECT	6.725 269.845 6.775 269.975 ;
		RECT	8.42 269.845 8.47 269.975 ;
		RECT	8.77 269.845 8.82 269.975 ;
		RECT	11.555 269.845 11.605 269.975 ;
		RECT	11.815 269.845 11.865 269.975 ;
		RECT	12.52 269.845 12.57 269.975 ;
		RECT	13.98 269.845 14.03 269.975 ;
		RECT	14.33 270.075 14.38 270.205 ;
		RECT	6.22 270.535 6.27 270.665 ;
		RECT	7.5 270.535 7.55 270.665 ;
		RECT	9.04 270.535 9.09 270.665 ;
		RECT	9.315 270.535 9.365 270.665 ;
		RECT	9.72 270.535 9.77 270.665 ;
		RECT	11.025 270.535 11.075 270.665 ;
		RECT	12.79 270.535 12.84 270.665 ;
		RECT	14.33 272.495 14.38 272.625 ;
		RECT	5.675 272.725 5.725 272.855 ;
		RECT	6.065 272.725 6.115 272.855 ;
		RECT	6.725 272.725 6.775 272.855 ;
		RECT	8.42 272.725 8.47 272.855 ;
		RECT	8.77 272.725 8.82 272.855 ;
		RECT	11.555 272.725 11.605 272.855 ;
		RECT	11.815 272.725 11.865 272.855 ;
		RECT	12.52 272.725 12.57 272.855 ;
		RECT	13.98 272.725 14.03 272.855 ;
		RECT	14.33 272.955 14.38 273.085 ;
		RECT	6.22 273.415 6.27 273.545 ;
		RECT	7.5 273.415 7.55 273.545 ;
		RECT	9.04 273.415 9.09 273.545 ;
		RECT	9.315 273.415 9.365 273.545 ;
		RECT	9.72 273.415 9.77 273.545 ;
		RECT	11.025 273.415 11.075 273.545 ;
		RECT	12.79 273.415 12.84 273.545 ;
		RECT	14.33 275.375 14.38 275.505 ;
		RECT	5.675 275.605 5.725 275.735 ;
		RECT	6.065 275.605 6.115 275.735 ;
		RECT	6.725 275.605 6.775 275.735 ;
		RECT	8.42 275.605 8.47 275.735 ;
		RECT	8.77 275.605 8.82 275.735 ;
		RECT	11.555 275.605 11.605 275.735 ;
		RECT	11.815 275.605 11.865 275.735 ;
		RECT	12.52 275.605 12.57 275.735 ;
		RECT	13.98 275.605 14.03 275.735 ;
		RECT	14.33 275.835 14.38 275.965 ;
		RECT	6.22 276.295 6.27 276.425 ;
		RECT	7.5 276.295 7.55 276.425 ;
		RECT	9.04 276.295 9.09 276.425 ;
		RECT	9.315 276.295 9.365 276.425 ;
		RECT	9.72 276.295 9.77 276.425 ;
		RECT	11.025 276.295 11.075 276.425 ;
		RECT	12.79 276.295 12.84 276.425 ;
		RECT	14.33 278.255 14.38 278.385 ;
		RECT	5.675 278.485 5.725 278.615 ;
		RECT	6.065 278.485 6.115 278.615 ;
		RECT	6.725 278.485 6.775 278.615 ;
		RECT	8.42 278.485 8.47 278.615 ;
		RECT	8.77 278.485 8.82 278.615 ;
		RECT	11.555 278.485 11.605 278.615 ;
		RECT	11.815 278.485 11.865 278.615 ;
		RECT	12.52 278.485 12.57 278.615 ;
		RECT	13.98 278.485 14.03 278.615 ;
		RECT	14.33 278.715 14.38 278.845 ;
		RECT	6.22 279.175 6.27 279.305 ;
		RECT	7.5 279.175 7.55 279.305 ;
		RECT	9.04 279.175 9.09 279.305 ;
		RECT	9.315 279.175 9.365 279.305 ;
		RECT	9.72 279.175 9.77 279.305 ;
		RECT	11.025 279.175 11.075 279.305 ;
		RECT	12.79 279.175 12.84 279.305 ;
		RECT	14.33 281.135 14.38 281.265 ;
		RECT	5.675 281.365 5.725 281.495 ;
		RECT	6.065 281.365 6.115 281.495 ;
		RECT	6.725 281.365 6.775 281.495 ;
		RECT	8.42 281.365 8.47 281.495 ;
		RECT	8.77 281.365 8.82 281.495 ;
		RECT	11.555 281.365 11.605 281.495 ;
		RECT	11.815 281.365 11.865 281.495 ;
		RECT	12.52 281.365 12.57 281.495 ;
		RECT	13.98 281.365 14.03 281.495 ;
		RECT	14.33 281.595 14.38 281.725 ;
		RECT	6.22 282.055 6.27 282.185 ;
		RECT	7.5 282.055 7.55 282.185 ;
		RECT	9.04 282.055 9.09 282.185 ;
		RECT	9.315 282.055 9.365 282.185 ;
		RECT	9.72 282.055 9.77 282.185 ;
		RECT	11.025 282.055 11.075 282.185 ;
		RECT	12.79 282.055 12.84 282.185 ;
		RECT	14.33 284.015 14.38 284.145 ;
		RECT	5.675 284.245 5.725 284.375 ;
		RECT	6.065 284.245 6.115 284.375 ;
		RECT	6.725 284.245 6.775 284.375 ;
		RECT	8.42 284.245 8.47 284.375 ;
		RECT	8.77 284.245 8.82 284.375 ;
		RECT	11.555 284.245 11.605 284.375 ;
		RECT	11.815 284.245 11.865 284.375 ;
		RECT	12.52 284.245 12.57 284.375 ;
		RECT	13.98 284.245 14.03 284.375 ;
		RECT	14.33 284.475 14.38 284.605 ;
		RECT	6.22 284.935 6.27 285.065 ;
		RECT	7.5 284.935 7.55 285.065 ;
		RECT	9.04 284.935 9.09 285.065 ;
		RECT	9.315 284.935 9.365 285.065 ;
		RECT	9.72 284.935 9.77 285.065 ;
		RECT	11.025 284.935 11.075 285.065 ;
		RECT	12.79 284.935 12.84 285.065 ;
		RECT	14.33 286.895 14.38 287.025 ;
		RECT	5.675 287.125 5.725 287.255 ;
		RECT	6.065 287.125 6.115 287.255 ;
		RECT	6.725 287.125 6.775 287.255 ;
		RECT	8.42 287.125 8.47 287.255 ;
		RECT	8.77 287.125 8.82 287.255 ;
		RECT	11.555 287.125 11.605 287.255 ;
		RECT	11.815 287.125 11.865 287.255 ;
		RECT	12.52 287.125 12.57 287.255 ;
		RECT	13.98 287.125 14.03 287.255 ;
		RECT	14.33 235.515 14.38 235.645 ;
		RECT	6.22 235.975 6.27 236.105 ;
		RECT	7.5 235.975 7.55 236.105 ;
		RECT	9.04 235.975 9.09 236.105 ;
		RECT	9.315 235.975 9.365 236.105 ;
		RECT	9.72 235.975 9.77 236.105 ;
		RECT	11.025 235.975 11.075 236.105 ;
		RECT	12.79 235.975 12.84 236.105 ;
		RECT	14.33 237.935 14.38 238.065 ;
		RECT	5.675 238.165 5.725 238.295 ;
		RECT	6.065 238.165 6.115 238.295 ;
		RECT	6.725 238.165 6.775 238.295 ;
		RECT	8.42 238.165 8.47 238.295 ;
		RECT	8.77 238.165 8.82 238.295 ;
		RECT	11.555 238.165 11.605 238.295 ;
		RECT	11.815 238.165 11.865 238.295 ;
		RECT	12.52 238.165 12.57 238.295 ;
		RECT	13.98 238.165 14.03 238.295 ;
		RECT	14.33 287.355 14.38 287.485 ;
		RECT	6.22 287.815 6.27 287.945 ;
		RECT	7.5 287.815 7.55 287.945 ;
		RECT	9.04 287.815 9.09 287.945 ;
		RECT	9.315 287.815 9.365 287.945 ;
		RECT	9.72 287.815 9.77 287.945 ;
		RECT	11.025 287.815 11.075 287.945 ;
		RECT	12.79 287.815 12.84 287.945 ;
		RECT	14.33 289.775 14.38 289.905 ;
		RECT	5.675 290.005 5.725 290.135 ;
		RECT	6.065 290.005 6.115 290.135 ;
		RECT	6.725 290.005 6.775 290.135 ;
		RECT	8.42 290.005 8.47 290.135 ;
		RECT	8.77 290.005 8.82 290.135 ;
		RECT	11.555 290.005 11.605 290.135 ;
		RECT	11.815 290.005 11.865 290.135 ;
		RECT	12.52 290.005 12.57 290.135 ;
		RECT	13.98 290.005 14.03 290.135 ;
		RECT	14.33 290.235 14.38 290.365 ;
		RECT	6.22 290.695 6.27 290.825 ;
		RECT	7.5 290.695 7.55 290.825 ;
		RECT	9.04 290.695 9.09 290.825 ;
		RECT	9.315 290.695 9.365 290.825 ;
		RECT	9.72 290.695 9.77 290.825 ;
		RECT	11.025 290.695 11.075 290.825 ;
		RECT	12.79 290.695 12.84 290.825 ;
		RECT	14.33 292.655 14.38 292.785 ;
		RECT	5.675 292.885 5.725 293.015 ;
		RECT	6.065 292.885 6.115 293.015 ;
		RECT	6.725 292.885 6.775 293.015 ;
		RECT	8.42 292.885 8.47 293.015 ;
		RECT	8.77 292.885 8.82 293.015 ;
		RECT	11.555 292.885 11.605 293.015 ;
		RECT	11.815 292.885 11.865 293.015 ;
		RECT	12.52 292.885 12.57 293.015 ;
		RECT	13.98 292.885 14.03 293.015 ;
		RECT	14.33 293.115 14.38 293.245 ;
		RECT	6.22 293.575 6.27 293.705 ;
		RECT	7.5 293.575 7.55 293.705 ;
		RECT	9.04 293.575 9.09 293.705 ;
		RECT	9.315 293.575 9.365 293.705 ;
		RECT	9.72 293.575 9.77 293.705 ;
		RECT	11.025 293.575 11.075 293.705 ;
		RECT	12.79 293.575 12.84 293.705 ;
		RECT	14.33 295.535 14.38 295.665 ;
		RECT	5.675 295.765 5.725 295.895 ;
		RECT	6.065 295.765 6.115 295.895 ;
		RECT	6.725 295.765 6.775 295.895 ;
		RECT	8.42 295.765 8.47 295.895 ;
		RECT	8.77 295.765 8.82 295.895 ;
		RECT	11.555 295.765 11.605 295.895 ;
		RECT	11.815 295.765 11.865 295.895 ;
		RECT	12.52 295.765 12.57 295.895 ;
		RECT	13.98 295.765 14.03 295.895 ;
		RECT	14.33 295.995 14.38 296.125 ;
		RECT	6.22 296.455 6.27 296.585 ;
		RECT	7.5 296.455 7.55 296.585 ;
		RECT	9.04 296.455 9.09 296.585 ;
		RECT	9.315 296.455 9.365 296.585 ;
		RECT	9.72 296.455 9.77 296.585 ;
		RECT	11.025 296.455 11.075 296.585 ;
		RECT	12.79 296.455 12.84 296.585 ;
		RECT	14.33 298.415 14.38 298.545 ;
		RECT	5.675 298.645 5.725 298.775 ;
		RECT	6.065 298.645 6.115 298.775 ;
		RECT	6.725 298.645 6.775 298.775 ;
		RECT	8.42 298.645 8.47 298.775 ;
		RECT	8.77 298.645 8.82 298.775 ;
		RECT	11.555 298.645 11.605 298.775 ;
		RECT	11.815 298.645 11.865 298.775 ;
		RECT	12.52 298.645 12.57 298.775 ;
		RECT	13.98 298.645 14.03 298.775 ;
		RECT	14.33 298.875 14.38 299.005 ;
		RECT	6.22 299.335 6.27 299.465 ;
		RECT	7.5 299.335 7.55 299.465 ;
		RECT	9.04 299.335 9.09 299.465 ;
		RECT	9.315 299.335 9.365 299.465 ;
		RECT	9.72 299.335 9.77 299.465 ;
		RECT	11.025 299.335 11.075 299.465 ;
		RECT	12.79 299.335 12.84 299.465 ;
		RECT	14.33 301.295 14.38 301.425 ;
		RECT	5.675 301.525 5.725 301.655 ;
		RECT	6.065 301.525 6.115 301.655 ;
		RECT	6.725 301.525 6.775 301.655 ;
		RECT	8.42 301.525 8.47 301.655 ;
		RECT	8.77 301.525 8.82 301.655 ;
		RECT	11.555 301.525 11.605 301.655 ;
		RECT	11.815 301.525 11.865 301.655 ;
		RECT	12.52 301.525 12.57 301.655 ;
		RECT	13.98 301.525 14.03 301.655 ;
		RECT	14.33 301.755 14.38 301.885 ;
		RECT	6.22 302.215 6.27 302.345 ;
		RECT	7.5 302.215 7.55 302.345 ;
		RECT	9.04 302.215 9.09 302.345 ;
		RECT	9.315 302.215 9.365 302.345 ;
		RECT	9.72 302.215 9.77 302.345 ;
		RECT	11.025 302.215 11.075 302.345 ;
		RECT	12.79 302.215 12.84 302.345 ;
		RECT	14.33 304.175 14.38 304.305 ;
		RECT	5.675 304.405 5.725 304.535 ;
		RECT	6.065 304.405 6.115 304.535 ;
		RECT	6.725 304.405 6.775 304.535 ;
		RECT	8.42 304.405 8.47 304.535 ;
		RECT	8.77 304.405 8.82 304.535 ;
		RECT	11.555 304.405 11.605 304.535 ;
		RECT	11.815 304.405 11.865 304.535 ;
		RECT	12.52 304.405 12.57 304.535 ;
		RECT	13.98 304.405 14.03 304.535 ;
		RECT	14.33 304.635 14.38 304.765 ;
		RECT	6.22 305.095 6.27 305.225 ;
		RECT	7.5 305.095 7.55 305.225 ;
		RECT	9.04 305.095 9.09 305.225 ;
		RECT	9.315 305.095 9.365 305.225 ;
		RECT	9.72 305.095 9.77 305.225 ;
		RECT	11.025 305.095 11.075 305.225 ;
		RECT	12.79 305.095 12.84 305.225 ;
		RECT	14.33 307.055 14.38 307.185 ;
		RECT	5.675 307.285 5.725 307.415 ;
		RECT	6.065 307.285 6.115 307.415 ;
		RECT	6.725 307.285 6.775 307.415 ;
		RECT	8.42 307.285 8.47 307.415 ;
		RECT	8.77 307.285 8.82 307.415 ;
		RECT	11.555 307.285 11.605 307.415 ;
		RECT	11.815 307.285 11.865 307.415 ;
		RECT	12.52 307.285 12.57 307.415 ;
		RECT	13.98 307.285 14.03 307.415 ;
		RECT	14.33 307.515 14.38 307.645 ;
		RECT	6.22 307.975 6.27 308.105 ;
		RECT	7.5 307.975 7.55 308.105 ;
		RECT	9.04 307.975 9.09 308.105 ;
		RECT	9.315 307.975 9.365 308.105 ;
		RECT	9.72 307.975 9.77 308.105 ;
		RECT	11.025 307.975 11.075 308.105 ;
		RECT	12.79 307.975 12.84 308.105 ;
		RECT	14.33 309.935 14.38 310.065 ;
		RECT	5.675 310.165 5.725 310.295 ;
		RECT	6.065 310.165 6.115 310.295 ;
		RECT	6.725 310.165 6.775 310.295 ;
		RECT	8.42 310.165 8.47 310.295 ;
		RECT	8.77 310.165 8.82 310.295 ;
		RECT	11.555 310.165 11.605 310.295 ;
		RECT	11.815 310.165 11.865 310.295 ;
		RECT	12.52 310.165 12.57 310.295 ;
		RECT	13.98 310.165 14.03 310.295 ;
		RECT	14.33 310.395 14.38 310.525 ;
		RECT	6.22 310.855 6.27 310.985 ;
		RECT	7.5 310.855 7.55 310.985 ;
		RECT	9.04 310.855 9.09 310.985 ;
		RECT	9.315 310.855 9.365 310.985 ;
		RECT	9.72 310.855 9.77 310.985 ;
		RECT	11.025 310.855 11.075 310.985 ;
		RECT	12.79 310.855 12.84 310.985 ;
		RECT	14.33 312.815 14.38 312.945 ;
		RECT	5.675 313.045 5.725 313.175 ;
		RECT	6.065 313.045 6.115 313.175 ;
		RECT	6.725 313.045 6.775 313.175 ;
		RECT	8.42 313.045 8.47 313.175 ;
		RECT	8.77 313.045 8.82 313.175 ;
		RECT	11.555 313.045 11.605 313.175 ;
		RECT	11.815 313.045 11.865 313.175 ;
		RECT	12.52 313.045 12.57 313.175 ;
		RECT	13.98 313.045 14.03 313.175 ;
		RECT	14.33 313.275 14.38 313.405 ;
		RECT	6.22 313.735 6.27 313.865 ;
		RECT	7.5 313.735 7.55 313.865 ;
		RECT	9.04 313.735 9.09 313.865 ;
		RECT	9.315 313.735 9.365 313.865 ;
		RECT	9.72 313.735 9.77 313.865 ;
		RECT	11.025 313.735 11.075 313.865 ;
		RECT	12.79 313.735 12.84 313.865 ;
		RECT	14.33 315.695 14.38 315.825 ;
		RECT	5.675 315.925 5.725 316.055 ;
		RECT	6.065 315.925 6.115 316.055 ;
		RECT	6.725 315.925 6.775 316.055 ;
		RECT	8.42 315.925 8.47 316.055 ;
		RECT	8.77 315.925 8.82 316.055 ;
		RECT	11.555 315.925 11.605 316.055 ;
		RECT	11.815 315.925 11.865 316.055 ;
		RECT	12.52 315.925 12.57 316.055 ;
		RECT	13.98 315.925 14.03 316.055 ;
		RECT	14.33 238.395 14.38 238.525 ;
		RECT	6.22 238.855 6.27 238.985 ;
		RECT	7.5 238.855 7.55 238.985 ;
		RECT	9.04 238.855 9.09 238.985 ;
		RECT	9.315 238.855 9.365 238.985 ;
		RECT	9.72 238.855 9.77 238.985 ;
		RECT	11.025 238.855 11.075 238.985 ;
		RECT	12.79 238.855 12.84 238.985 ;
		RECT	14.33 240.815 14.38 240.945 ;
		RECT	5.675 241.045 5.725 241.175 ;
		RECT	6.065 241.045 6.115 241.175 ;
		RECT	6.725 241.045 6.775 241.175 ;
		RECT	8.42 241.045 8.47 241.175 ;
		RECT	8.77 241.045 8.82 241.175 ;
		RECT	11.555 241.045 11.605 241.175 ;
		RECT	11.815 241.045 11.865 241.175 ;
		RECT	12.52 241.045 12.57 241.175 ;
		RECT	13.98 241.045 14.03 241.175 ;
		RECT	14.33 316.155 14.38 316.285 ;
		RECT	6.22 316.615 6.27 316.745 ;
		RECT	7.5 316.615 7.55 316.745 ;
		RECT	9.04 316.615 9.09 316.745 ;
		RECT	9.315 316.615 9.365 316.745 ;
		RECT	9.72 316.615 9.77 316.745 ;
		RECT	11.025 316.615 11.075 316.745 ;
		RECT	12.79 316.615 12.84 316.745 ;
		RECT	14.33 318.575 14.38 318.705 ;
		RECT	5.675 318.805 5.725 318.935 ;
		RECT	6.065 318.805 6.115 318.935 ;
		RECT	6.725 318.805 6.775 318.935 ;
		RECT	8.42 318.805 8.47 318.935 ;
		RECT	8.77 318.805 8.82 318.935 ;
		RECT	11.555 318.805 11.605 318.935 ;
		RECT	11.815 318.805 11.865 318.935 ;
		RECT	12.52 318.805 12.57 318.935 ;
		RECT	13.98 318.805 14.03 318.935 ;
		RECT	14.33 319.035 14.38 319.165 ;
		RECT	6.22 319.495 6.27 319.625 ;
		RECT	7.5 319.495 7.55 319.625 ;
		RECT	9.04 319.495 9.09 319.625 ;
		RECT	9.315 319.495 9.365 319.625 ;
		RECT	9.72 319.495 9.77 319.625 ;
		RECT	11.025 319.495 11.075 319.625 ;
		RECT	12.79 319.495 12.84 319.625 ;
		RECT	14.33 321.455 14.38 321.585 ;
		RECT	5.675 321.685 5.725 321.815 ;
		RECT	6.065 321.685 6.115 321.815 ;
		RECT	6.725 321.685 6.775 321.815 ;
		RECT	8.42 321.685 8.47 321.815 ;
		RECT	8.77 321.685 8.82 321.815 ;
		RECT	11.555 321.685 11.605 321.815 ;
		RECT	11.815 321.685 11.865 321.815 ;
		RECT	12.52 321.685 12.57 321.815 ;
		RECT	13.98 321.685 14.03 321.815 ;
		RECT	14.33 321.915 14.38 322.045 ;
		RECT	6.22 322.375 6.27 322.505 ;
		RECT	7.5 322.375 7.55 322.505 ;
		RECT	9.04 322.375 9.09 322.505 ;
		RECT	9.315 322.375 9.365 322.505 ;
		RECT	9.72 322.375 9.77 322.505 ;
		RECT	11.025 322.375 11.075 322.505 ;
		RECT	12.79 322.375 12.84 322.505 ;
		RECT	14.33 324.335 14.38 324.465 ;
		RECT	5.675 324.565 5.725 324.695 ;
		RECT	6.065 324.565 6.115 324.695 ;
		RECT	6.725 324.565 6.775 324.695 ;
		RECT	8.42 324.565 8.47 324.695 ;
		RECT	8.77 324.565 8.82 324.695 ;
		RECT	11.555 324.565 11.605 324.695 ;
		RECT	11.815 324.565 11.865 324.695 ;
		RECT	12.52 324.565 12.57 324.695 ;
		RECT	13.98 324.565 14.03 324.695 ;
		RECT	14.33 324.795 14.38 324.925 ;
		RECT	6.22 325.255 6.27 325.385 ;
		RECT	7.5 325.255 7.55 325.385 ;
		RECT	9.04 325.255 9.09 325.385 ;
		RECT	9.315 325.255 9.365 325.385 ;
		RECT	9.72 325.255 9.77 325.385 ;
		RECT	11.025 325.255 11.075 325.385 ;
		RECT	12.79 325.255 12.84 325.385 ;
		RECT	14.33 327.215 14.38 327.345 ;
		RECT	5.675 327.445 5.725 327.575 ;
		RECT	6.065 327.445 6.115 327.575 ;
		RECT	6.725 327.445 6.775 327.575 ;
		RECT	8.42 327.445 8.47 327.575 ;
		RECT	8.77 327.445 8.82 327.575 ;
		RECT	11.555 327.445 11.605 327.575 ;
		RECT	11.815 327.445 11.865 327.575 ;
		RECT	12.52 327.445 12.57 327.575 ;
		RECT	13.98 327.445 14.03 327.575 ;
		RECT	14.33 327.675 14.38 327.805 ;
		RECT	6.22 328.135 6.27 328.265 ;
		RECT	7.5 328.135 7.55 328.265 ;
		RECT	9.04 328.135 9.09 328.265 ;
		RECT	9.315 328.135 9.365 328.265 ;
		RECT	9.72 328.135 9.77 328.265 ;
		RECT	11.025 328.135 11.075 328.265 ;
		RECT	12.79 328.135 12.84 328.265 ;
		RECT	14.33 330.095 14.38 330.225 ;
		RECT	5.675 330.325 5.725 330.455 ;
		RECT	6.065 330.325 6.115 330.455 ;
		RECT	6.725 330.325 6.775 330.455 ;
		RECT	8.42 330.325 8.47 330.455 ;
		RECT	8.77 330.325 8.82 330.455 ;
		RECT	11.555 330.325 11.605 330.455 ;
		RECT	11.815 330.325 11.865 330.455 ;
		RECT	12.52 330.325 12.57 330.455 ;
		RECT	13.98 330.325 14.03 330.455 ;
		RECT	14.33 330.555 14.38 330.685 ;
		RECT	6.22 331.015 6.27 331.145 ;
		RECT	7.5 331.015 7.55 331.145 ;
		RECT	9.04 331.015 9.09 331.145 ;
		RECT	9.315 331.015 9.365 331.145 ;
		RECT	9.72 331.015 9.77 331.145 ;
		RECT	11.025 331.015 11.075 331.145 ;
		RECT	12.79 331.015 12.84 331.145 ;
		RECT	14.33 332.975 14.38 333.105 ;
		RECT	5.675 333.205 5.725 333.335 ;
		RECT	6.065 333.205 6.115 333.335 ;
		RECT	6.725 333.205 6.775 333.335 ;
		RECT	8.42 333.205 8.47 333.335 ;
		RECT	8.77 333.205 8.82 333.335 ;
		RECT	11.555 333.205 11.605 333.335 ;
		RECT	11.815 333.205 11.865 333.335 ;
		RECT	12.52 333.205 12.57 333.335 ;
		RECT	13.98 333.205 14.03 333.335 ;
		RECT	14.33 333.435 14.38 333.565 ;
		RECT	6.22 333.895 6.27 334.025 ;
		RECT	7.5 333.895 7.55 334.025 ;
		RECT	9.04 333.895 9.09 334.025 ;
		RECT	9.315 333.895 9.365 334.025 ;
		RECT	9.72 333.895 9.77 334.025 ;
		RECT	11.025 333.895 11.075 334.025 ;
		RECT	12.79 333.895 12.84 334.025 ;
		RECT	14.33 335.855 14.38 335.985 ;
		RECT	5.675 336.085 5.725 336.215 ;
		RECT	6.065 336.085 6.115 336.215 ;
		RECT	6.725 336.085 6.775 336.215 ;
		RECT	8.42 336.085 8.47 336.215 ;
		RECT	8.77 336.085 8.82 336.215 ;
		RECT	11.555 336.085 11.605 336.215 ;
		RECT	11.815 336.085 11.865 336.215 ;
		RECT	12.52 336.085 12.57 336.215 ;
		RECT	13.98 336.085 14.03 336.215 ;
		RECT	14.33 336.315 14.38 336.445 ;
		RECT	6.22 336.775 6.27 336.905 ;
		RECT	7.5 336.775 7.55 336.905 ;
		RECT	9.04 336.775 9.09 336.905 ;
		RECT	9.315 336.775 9.365 336.905 ;
		RECT	9.72 336.775 9.77 336.905 ;
		RECT	11.025 336.775 11.075 336.905 ;
		RECT	12.79 336.775 12.84 336.905 ;
		RECT	14.33 338.735 14.38 338.865 ;
		RECT	5.675 338.965 5.725 339.095 ;
		RECT	6.065 338.965 6.115 339.095 ;
		RECT	6.725 338.965 6.775 339.095 ;
		RECT	8.42 338.965 8.47 339.095 ;
		RECT	8.77 338.965 8.82 339.095 ;
		RECT	11.555 338.965 11.605 339.095 ;
		RECT	11.815 338.965 11.865 339.095 ;
		RECT	12.52 338.965 12.57 339.095 ;
		RECT	13.98 338.965 14.03 339.095 ;
		RECT	14.33 339.195 14.38 339.325 ;
		RECT	6.22 339.655 6.27 339.785 ;
		RECT	7.5 339.655 7.55 339.785 ;
		RECT	9.04 339.655 9.09 339.785 ;
		RECT	9.315 339.655 9.365 339.785 ;
		RECT	9.72 339.655 9.77 339.785 ;
		RECT	11.025 339.655 11.075 339.785 ;
		RECT	12.79 339.655 12.84 339.785 ;
		RECT	14.33 341.615 14.38 341.745 ;
		RECT	5.675 341.845 5.725 341.975 ;
		RECT	6.065 341.845 6.115 341.975 ;
		RECT	6.725 341.845 6.775 341.975 ;
		RECT	8.42 341.845 8.47 341.975 ;
		RECT	8.77 341.845 8.82 341.975 ;
		RECT	11.555 341.845 11.605 341.975 ;
		RECT	11.815 341.845 11.865 341.975 ;
		RECT	12.52 341.845 12.57 341.975 ;
		RECT	13.98 341.845 14.03 341.975 ;
		RECT	14.33 342.075 14.38 342.205 ;
		RECT	6.22 342.535 6.27 342.665 ;
		RECT	7.5 342.535 7.55 342.665 ;
		RECT	9.04 342.535 9.09 342.665 ;
		RECT	9.315 342.535 9.365 342.665 ;
		RECT	9.72 342.535 9.77 342.665 ;
		RECT	11.025 342.535 11.075 342.665 ;
		RECT	12.79 342.535 12.84 342.665 ;
		RECT	14.33 344.495 14.38 344.625 ;
		RECT	5.675 344.725 5.725 344.855 ;
		RECT	6.065 344.725 6.115 344.855 ;
		RECT	6.725 344.725 6.775 344.855 ;
		RECT	8.42 344.725 8.47 344.855 ;
		RECT	8.77 344.725 8.82 344.855 ;
		RECT	11.555 344.725 11.605 344.855 ;
		RECT	11.815 344.725 11.865 344.855 ;
		RECT	12.52 344.725 12.57 344.855 ;
		RECT	13.98 344.725 14.03 344.855 ;
		RECT	14.33 241.275 14.38 241.405 ;
		RECT	6.22 241.735 6.27 241.865 ;
		RECT	7.5 241.735 7.55 241.865 ;
		RECT	9.04 241.735 9.09 241.865 ;
		RECT	9.315 241.735 9.365 241.865 ;
		RECT	9.72 241.735 9.77 241.865 ;
		RECT	11.025 241.735 11.075 241.865 ;
		RECT	12.79 241.735 12.84 241.865 ;
		RECT	14.33 243.695 14.38 243.825 ;
		RECT	5.675 243.925 5.725 244.055 ;
		RECT	6.065 243.925 6.115 244.055 ;
		RECT	6.725 243.925 6.775 244.055 ;
		RECT	8.42 243.925 8.47 244.055 ;
		RECT	8.77 243.925 8.82 244.055 ;
		RECT	11.555 243.925 11.605 244.055 ;
		RECT	11.815 243.925 11.865 244.055 ;
		RECT	12.52 243.925 12.57 244.055 ;
		RECT	13.98 243.925 14.03 244.055 ;
		RECT	14.33 344.955 14.38 345.085 ;
		RECT	6.22 345.415 6.27 345.545 ;
		RECT	7.5 345.415 7.55 345.545 ;
		RECT	9.04 345.415 9.09 345.545 ;
		RECT	9.315 345.415 9.365 345.545 ;
		RECT	9.72 345.415 9.77 345.545 ;
		RECT	11.025 345.415 11.075 345.545 ;
		RECT	12.79 345.415 12.84 345.545 ;
		RECT	14.33 347.375 14.38 347.505 ;
		RECT	5.675 347.605 5.725 347.735 ;
		RECT	6.065 347.605 6.115 347.735 ;
		RECT	6.725 347.605 6.775 347.735 ;
		RECT	8.42 347.605 8.47 347.735 ;
		RECT	8.77 347.605 8.82 347.735 ;
		RECT	11.555 347.605 11.605 347.735 ;
		RECT	11.815 347.605 11.865 347.735 ;
		RECT	12.52 347.605 12.57 347.735 ;
		RECT	13.98 347.605 14.03 347.735 ;
		RECT	14.33 347.835 14.38 347.965 ;
		RECT	6.22 348.295 6.27 348.425 ;
		RECT	7.5 348.295 7.55 348.425 ;
		RECT	9.04 348.295 9.09 348.425 ;
		RECT	9.315 348.295 9.365 348.425 ;
		RECT	9.72 348.295 9.77 348.425 ;
		RECT	11.025 348.295 11.075 348.425 ;
		RECT	12.79 348.295 12.84 348.425 ;
		RECT	14.33 350.255 14.38 350.385 ;
		RECT	5.675 350.485 5.725 350.615 ;
		RECT	6.065 350.485 6.115 350.615 ;
		RECT	6.725 350.485 6.775 350.615 ;
		RECT	8.42 350.485 8.47 350.615 ;
		RECT	8.77 350.485 8.82 350.615 ;
		RECT	11.555 350.485 11.605 350.615 ;
		RECT	11.815 350.485 11.865 350.615 ;
		RECT	12.52 350.485 12.57 350.615 ;
		RECT	13.98 350.485 14.03 350.615 ;
		RECT	14.33 350.715 14.38 350.845 ;
		RECT	6.22 351.175 6.27 351.305 ;
		RECT	7.5 351.175 7.55 351.305 ;
		RECT	9.04 351.175 9.09 351.305 ;
		RECT	9.315 351.175 9.365 351.305 ;
		RECT	9.72 351.175 9.77 351.305 ;
		RECT	11.025 351.175 11.075 351.305 ;
		RECT	12.79 351.175 12.84 351.305 ;
		RECT	14.33 353.135 14.38 353.265 ;
		RECT	5.675 353.365 5.725 353.495 ;
		RECT	6.065 353.365 6.115 353.495 ;
		RECT	6.725 353.365 6.775 353.495 ;
		RECT	8.42 353.365 8.47 353.495 ;
		RECT	8.77 353.365 8.82 353.495 ;
		RECT	11.555 353.365 11.605 353.495 ;
		RECT	11.815 353.365 11.865 353.495 ;
		RECT	12.52 353.365 12.57 353.495 ;
		RECT	13.98 353.365 14.03 353.495 ;
		RECT	14.33 353.595 14.38 353.725 ;
		RECT	6.22 354.055 6.27 354.185 ;
		RECT	7.5 354.055 7.55 354.185 ;
		RECT	9.04 354.055 9.09 354.185 ;
		RECT	9.315 354.055 9.365 354.185 ;
		RECT	9.72 354.055 9.77 354.185 ;
		RECT	11.025 354.055 11.075 354.185 ;
		RECT	12.79 354.055 12.84 354.185 ;
		RECT	14.33 356.015 14.38 356.145 ;
		RECT	5.675 356.245 5.725 356.375 ;
		RECT	6.065 356.245 6.115 356.375 ;
		RECT	6.725 356.245 6.775 356.375 ;
		RECT	8.42 356.245 8.47 356.375 ;
		RECT	8.77 356.245 8.82 356.375 ;
		RECT	11.555 356.245 11.605 356.375 ;
		RECT	11.815 356.245 11.865 356.375 ;
		RECT	12.52 356.245 12.57 356.375 ;
		RECT	13.98 356.245 14.03 356.375 ;
		RECT	14.33 356.475 14.38 356.605 ;
		RECT	6.22 356.935 6.27 357.065 ;
		RECT	7.5 356.935 7.55 357.065 ;
		RECT	9.04 356.935 9.09 357.065 ;
		RECT	9.315 356.935 9.365 357.065 ;
		RECT	9.72 356.935 9.77 357.065 ;
		RECT	11.025 356.935 11.075 357.065 ;
		RECT	12.79 356.935 12.84 357.065 ;
		RECT	14.33 358.895 14.38 359.025 ;
		RECT	5.675 359.125 5.725 359.255 ;
		RECT	6.065 359.125 6.115 359.255 ;
		RECT	6.725 359.125 6.775 359.255 ;
		RECT	8.42 359.125 8.47 359.255 ;
		RECT	8.77 359.125 8.82 359.255 ;
		RECT	11.555 359.125 11.605 359.255 ;
		RECT	11.815 359.125 11.865 359.255 ;
		RECT	12.52 359.125 12.57 359.255 ;
		RECT	13.98 359.125 14.03 359.255 ;
		RECT	14.33 359.355 14.38 359.485 ;
		RECT	6.22 359.815 6.27 359.945 ;
		RECT	7.5 359.815 7.55 359.945 ;
		RECT	9.04 359.815 9.09 359.945 ;
		RECT	9.315 359.815 9.365 359.945 ;
		RECT	9.72 359.815 9.77 359.945 ;
		RECT	11.025 359.815 11.075 359.945 ;
		RECT	12.79 359.815 12.84 359.945 ;
		RECT	14.33 361.775 14.38 361.905 ;
		RECT	5.675 362.005 5.725 362.135 ;
		RECT	6.065 362.005 6.115 362.135 ;
		RECT	6.725 362.005 6.775 362.135 ;
		RECT	8.42 362.005 8.47 362.135 ;
		RECT	8.77 362.005 8.82 362.135 ;
		RECT	11.555 362.005 11.605 362.135 ;
		RECT	11.815 362.005 11.865 362.135 ;
		RECT	12.52 362.005 12.57 362.135 ;
		RECT	13.98 362.005 14.03 362.135 ;
		RECT	14.33 362.235 14.38 362.365 ;
		RECT	6.22 362.695 6.27 362.825 ;
		RECT	7.5 362.695 7.55 362.825 ;
		RECT	9.04 362.695 9.09 362.825 ;
		RECT	9.315 362.695 9.365 362.825 ;
		RECT	9.72 362.695 9.77 362.825 ;
		RECT	11.025 362.695 11.075 362.825 ;
		RECT	12.79 362.695 12.84 362.825 ;
		RECT	14.33 364.655 14.38 364.785 ;
		RECT	5.675 364.885 5.725 365.015 ;
		RECT	6.065 364.885 6.115 365.015 ;
		RECT	6.725 364.885 6.775 365.015 ;
		RECT	8.42 364.885 8.47 365.015 ;
		RECT	8.77 364.885 8.82 365.015 ;
		RECT	11.555 364.885 11.605 365.015 ;
		RECT	11.815 364.885 11.865 365.015 ;
		RECT	12.52 364.885 12.57 365.015 ;
		RECT	13.98 364.885 14.03 365.015 ;
		RECT	14.33 365.115 14.38 365.245 ;
		RECT	6.22 365.575 6.27 365.705 ;
		RECT	7.5 365.575 7.55 365.705 ;
		RECT	9.04 365.575 9.09 365.705 ;
		RECT	9.315 365.575 9.365 365.705 ;
		RECT	9.72 365.575 9.77 365.705 ;
		RECT	11.025 365.575 11.075 365.705 ;
		RECT	12.79 365.575 12.84 365.705 ;
		RECT	14.33 367.535 14.38 367.665 ;
		RECT	5.675 367.765 5.725 367.895 ;
		RECT	6.065 367.765 6.115 367.895 ;
		RECT	6.725 367.765 6.775 367.895 ;
		RECT	8.42 367.765 8.47 367.895 ;
		RECT	8.77 367.765 8.82 367.895 ;
		RECT	11.555 367.765 11.605 367.895 ;
		RECT	11.815 367.765 11.865 367.895 ;
		RECT	12.52 367.765 12.57 367.895 ;
		RECT	13.98 367.765 14.03 367.895 ;
		RECT	14.33 367.995 14.38 368.125 ;
		RECT	6.22 368.455 6.27 368.585 ;
		RECT	7.5 368.455 7.55 368.585 ;
		RECT	9.04 368.455 9.09 368.585 ;
		RECT	9.315 368.455 9.365 368.585 ;
		RECT	9.72 368.455 9.77 368.585 ;
		RECT	11.025 368.455 11.075 368.585 ;
		RECT	12.79 368.455 12.84 368.585 ;
		RECT	14.33 370.415 14.38 370.545 ;
		RECT	5.675 370.645 5.725 370.775 ;
		RECT	6.065 370.645 6.115 370.775 ;
		RECT	6.725 370.645 6.775 370.775 ;
		RECT	8.42 370.645 8.47 370.775 ;
		RECT	8.77 370.645 8.82 370.775 ;
		RECT	11.555 370.645 11.605 370.775 ;
		RECT	11.815 370.645 11.865 370.775 ;
		RECT	12.52 370.645 12.57 370.775 ;
		RECT	13.98 370.645 14.03 370.775 ;
		RECT	14.33 370.875 14.38 371.005 ;
		RECT	6.22 371.335 6.27 371.465 ;
		RECT	7.5 371.335 7.55 371.465 ;
		RECT	9.04 371.335 9.09 371.465 ;
		RECT	9.315 371.335 9.365 371.465 ;
		RECT	9.72 371.335 9.77 371.465 ;
		RECT	11.025 371.335 11.075 371.465 ;
		RECT	12.79 371.335 12.84 371.465 ;
		RECT	14.33 373.295 14.38 373.425 ;
		RECT	5.675 373.525 5.725 373.655 ;
		RECT	6.065 373.525 6.115 373.655 ;
		RECT	6.725 373.525 6.775 373.655 ;
		RECT	8.42 373.525 8.47 373.655 ;
		RECT	8.77 373.525 8.82 373.655 ;
		RECT	11.555 373.525 11.605 373.655 ;
		RECT	11.815 373.525 11.865 373.655 ;
		RECT	12.52 373.525 12.57 373.655 ;
		RECT	13.98 373.525 14.03 373.655 ;
		RECT	14.33 244.155 14.38 244.285 ;
		RECT	6.22 244.615 6.27 244.745 ;
		RECT	7.5 244.615 7.55 244.745 ;
		RECT	9.04 244.615 9.09 244.745 ;
		RECT	9.315 244.615 9.365 244.745 ;
		RECT	9.72 244.615 9.77 244.745 ;
		RECT	11.025 244.615 11.075 244.745 ;
		RECT	12.79 244.615 12.84 244.745 ;
		RECT	14.33 246.575 14.38 246.705 ;
		RECT	5.675 246.805 5.725 246.935 ;
		RECT	6.065 246.805 6.115 246.935 ;
		RECT	6.725 246.805 6.775 246.935 ;
		RECT	8.42 246.805 8.47 246.935 ;
		RECT	8.77 246.805 8.82 246.935 ;
		RECT	11.555 246.805 11.605 246.935 ;
		RECT	11.815 246.805 11.865 246.935 ;
		RECT	12.52 246.805 12.57 246.935 ;
		RECT	13.98 246.805 14.03 246.935 ;
		RECT	14.33 373.755 14.38 373.885 ;
		RECT	6.22 374.215 6.27 374.345 ;
		RECT	7.5 374.215 7.55 374.345 ;
		RECT	9.04 374.215 9.09 374.345 ;
		RECT	9.315 374.215 9.365 374.345 ;
		RECT	9.72 374.215 9.77 374.345 ;
		RECT	11.025 374.215 11.075 374.345 ;
		RECT	12.79 374.215 12.84 374.345 ;
		RECT	14.33 376.175 14.38 376.305 ;
		RECT	5.675 376.405 5.725 376.535 ;
		RECT	6.065 376.405 6.115 376.535 ;
		RECT	6.725 376.405 6.775 376.535 ;
		RECT	8.42 376.405 8.47 376.535 ;
		RECT	8.77 376.405 8.82 376.535 ;
		RECT	11.555 376.405 11.605 376.535 ;
		RECT	11.815 376.405 11.865 376.535 ;
		RECT	12.52 376.405 12.57 376.535 ;
		RECT	13.98 376.405 14.03 376.535 ;
		RECT	14.33 376.635 14.38 376.765 ;
		RECT	6.22 377.095 6.27 377.225 ;
		RECT	7.5 377.095 7.55 377.225 ;
		RECT	9.04 377.095 9.09 377.225 ;
		RECT	9.315 377.095 9.365 377.225 ;
		RECT	9.72 377.095 9.77 377.225 ;
		RECT	11.025 377.095 11.075 377.225 ;
		RECT	12.79 377.095 12.84 377.225 ;
		RECT	14.33 379.055 14.38 379.185 ;
		RECT	5.675 379.285 5.725 379.415 ;
		RECT	6.065 379.285 6.115 379.415 ;
		RECT	6.725 379.285 6.775 379.415 ;
		RECT	8.42 379.285 8.47 379.415 ;
		RECT	8.77 379.285 8.82 379.415 ;
		RECT	11.555 379.285 11.605 379.415 ;
		RECT	11.815 379.285 11.865 379.415 ;
		RECT	12.52 379.285 12.57 379.415 ;
		RECT	13.98 379.285 14.03 379.415 ;
		RECT	14.33 379.515 14.38 379.645 ;
		RECT	6.22 379.975 6.27 380.105 ;
		RECT	7.5 379.975 7.55 380.105 ;
		RECT	9.04 379.975 9.09 380.105 ;
		RECT	9.315 379.975 9.365 380.105 ;
		RECT	9.72 379.975 9.77 380.105 ;
		RECT	11.025 379.975 11.075 380.105 ;
		RECT	12.79 379.975 12.84 380.105 ;
		RECT	14.33 381.935 14.38 382.065 ;
		RECT	5.675 382.165 5.725 382.295 ;
		RECT	6.065 382.165 6.115 382.295 ;
		RECT	6.725 382.165 6.775 382.295 ;
		RECT	8.42 382.165 8.47 382.295 ;
		RECT	8.77 382.165 8.82 382.295 ;
		RECT	11.555 382.165 11.605 382.295 ;
		RECT	11.815 382.165 11.865 382.295 ;
		RECT	12.52 382.165 12.57 382.295 ;
		RECT	13.98 382.165 14.03 382.295 ;
		RECT	14.33 382.395 14.38 382.525 ;
		RECT	6.22 382.855 6.27 382.985 ;
		RECT	7.5 382.855 7.55 382.985 ;
		RECT	9.04 382.855 9.09 382.985 ;
		RECT	9.315 382.855 9.365 382.985 ;
		RECT	9.72 382.855 9.77 382.985 ;
		RECT	11.025 382.855 11.075 382.985 ;
		RECT	12.79 382.855 12.84 382.985 ;
		RECT	14.33 384.815 14.38 384.945 ;
		RECT	5.675 385.045 5.725 385.175 ;
		RECT	6.065 385.045 6.115 385.175 ;
		RECT	6.725 385.045 6.775 385.175 ;
		RECT	8.42 385.045 8.47 385.175 ;
		RECT	8.77 385.045 8.82 385.175 ;
		RECT	11.555 385.045 11.605 385.175 ;
		RECT	11.815 385.045 11.865 385.175 ;
		RECT	12.52 385.045 12.57 385.175 ;
		RECT	13.98 385.045 14.03 385.175 ;
		RECT	14.33 385.275 14.38 385.405 ;
		RECT	6.22 385.735 6.27 385.865 ;
		RECT	7.5 385.735 7.55 385.865 ;
		RECT	9.04 385.735 9.09 385.865 ;
		RECT	9.315 385.735 9.365 385.865 ;
		RECT	9.72 385.735 9.77 385.865 ;
		RECT	11.025 385.735 11.075 385.865 ;
		RECT	12.79 385.735 12.84 385.865 ;
		RECT	14.33 387.695 14.38 387.825 ;
		RECT	5.675 387.925 5.725 388.055 ;
		RECT	6.065 387.925 6.115 388.055 ;
		RECT	6.725 387.925 6.775 388.055 ;
		RECT	8.42 387.925 8.47 388.055 ;
		RECT	8.77 387.925 8.82 388.055 ;
		RECT	11.555 387.925 11.605 388.055 ;
		RECT	11.815 387.925 11.865 388.055 ;
		RECT	12.52 387.925 12.57 388.055 ;
		RECT	13.98 387.925 14.03 388.055 ;
		RECT	14.33 388.155 14.38 388.285 ;
		RECT	6.22 388.615 6.27 388.745 ;
		RECT	7.5 388.615 7.55 388.745 ;
		RECT	9.04 388.615 9.09 388.745 ;
		RECT	9.315 388.615 9.365 388.745 ;
		RECT	9.72 388.615 9.77 388.745 ;
		RECT	11.025 388.615 11.075 388.745 ;
		RECT	12.79 388.615 12.84 388.745 ;
		RECT	14.33 390.575 14.38 390.705 ;
		RECT	5.675 390.805 5.725 390.935 ;
		RECT	6.065 390.805 6.115 390.935 ;
		RECT	6.725 390.805 6.775 390.935 ;
		RECT	8.42 390.805 8.47 390.935 ;
		RECT	8.77 390.805 8.82 390.935 ;
		RECT	11.555 390.805 11.605 390.935 ;
		RECT	11.815 390.805 11.865 390.935 ;
		RECT	12.52 390.805 12.57 390.935 ;
		RECT	13.98 390.805 14.03 390.935 ;
		RECT	14.33 391.035 14.38 391.165 ;
		RECT	6.22 391.495 6.27 391.625 ;
		RECT	7.5 391.495 7.55 391.625 ;
		RECT	9.04 391.495 9.09 391.625 ;
		RECT	9.315 391.495 9.365 391.625 ;
		RECT	9.72 391.495 9.77 391.625 ;
		RECT	11.025 391.495 11.075 391.625 ;
		RECT	12.79 391.495 12.84 391.625 ;
		RECT	14.33 393.455 14.38 393.585 ;
		RECT	5.675 393.685 5.725 393.815 ;
		RECT	6.065 393.685 6.115 393.815 ;
		RECT	6.725 393.685 6.775 393.815 ;
		RECT	8.42 393.685 8.47 393.815 ;
		RECT	8.77 393.685 8.82 393.815 ;
		RECT	11.555 393.685 11.605 393.815 ;
		RECT	11.815 393.685 11.865 393.815 ;
		RECT	12.52 393.685 12.57 393.815 ;
		RECT	13.98 393.685 14.03 393.815 ;
		RECT	14.33 393.915 14.38 394.045 ;
		RECT	6.22 394.375 6.27 394.505 ;
		RECT	7.5 394.375 7.55 394.505 ;
		RECT	9.04 394.375 9.09 394.505 ;
		RECT	9.315 394.375 9.365 394.505 ;
		RECT	9.72 394.375 9.77 394.505 ;
		RECT	11.025 394.375 11.075 394.505 ;
		RECT	12.79 394.375 12.84 394.505 ;
		RECT	14.33 396.335 14.38 396.465 ;
		RECT	5.675 396.565 5.725 396.695 ;
		RECT	6.065 396.565 6.115 396.695 ;
		RECT	6.725 396.565 6.775 396.695 ;
		RECT	8.42 396.565 8.47 396.695 ;
		RECT	8.77 396.565 8.82 396.695 ;
		RECT	11.555 396.565 11.605 396.695 ;
		RECT	11.815 396.565 11.865 396.695 ;
		RECT	12.52 396.565 12.57 396.695 ;
		RECT	13.98 396.565 14.03 396.695 ;
		RECT	14.33 396.795 14.38 396.925 ;
		RECT	6.22 397.255 6.27 397.385 ;
		RECT	7.5 397.255 7.55 397.385 ;
		RECT	9.04 397.255 9.09 397.385 ;
		RECT	9.315 397.255 9.365 397.385 ;
		RECT	9.72 397.255 9.77 397.385 ;
		RECT	11.025 397.255 11.075 397.385 ;
		RECT	12.79 397.255 12.84 397.385 ;
		RECT	14.33 399.215 14.38 399.345 ;
		RECT	5.675 399.445 5.725 399.575 ;
		RECT	6.065 399.445 6.115 399.575 ;
		RECT	6.725 399.445 6.775 399.575 ;
		RECT	8.42 399.445 8.47 399.575 ;
		RECT	8.77 399.445 8.82 399.575 ;
		RECT	11.555 399.445 11.605 399.575 ;
		RECT	11.815 399.445 11.865 399.575 ;
		RECT	12.52 399.445 12.57 399.575 ;
		RECT	13.98 399.445 14.03 399.575 ;
		RECT	14.33 399.675 14.38 399.805 ;
		RECT	6.22 400.135 6.27 400.265 ;
		RECT	7.5 400.135 7.55 400.265 ;
		RECT	9.04 400.135 9.09 400.265 ;
		RECT	9.315 400.135 9.365 400.265 ;
		RECT	9.72 400.135 9.77 400.265 ;
		RECT	11.025 400.135 11.075 400.265 ;
		RECT	12.79 400.135 12.84 400.265 ;
		RECT	14.33 402.095 14.38 402.225 ;
		RECT	5.675 402.325 5.725 402.455 ;
		RECT	6.065 402.325 6.115 402.455 ;
		RECT	6.725 402.325 6.775 402.455 ;
		RECT	8.42 402.325 8.47 402.455 ;
		RECT	8.77 402.325 8.82 402.455 ;
		RECT	11.555 402.325 11.605 402.455 ;
		RECT	11.815 402.325 11.865 402.455 ;
		RECT	12.52 402.325 12.57 402.455 ;
		RECT	13.98 402.325 14.03 402.455 ;
		RECT	14.33 247.035 14.38 247.165 ;
		RECT	6.22 247.495 6.27 247.625 ;
		RECT	7.5 247.495 7.55 247.625 ;
		RECT	9.04 247.495 9.09 247.625 ;
		RECT	9.315 247.495 9.365 247.625 ;
		RECT	9.72 247.495 9.77 247.625 ;
		RECT	11.025 247.495 11.075 247.625 ;
		RECT	12.79 247.495 12.84 247.625 ;
		RECT	14.33 249.455 14.38 249.585 ;
		RECT	5.675 249.685 5.725 249.815 ;
		RECT	6.065 249.685 6.115 249.815 ;
		RECT	6.725 249.685 6.775 249.815 ;
		RECT	8.42 249.685 8.47 249.815 ;
		RECT	8.77 249.685 8.82 249.815 ;
		RECT	11.555 249.685 11.605 249.815 ;
		RECT	11.815 249.685 11.865 249.815 ;
		RECT	12.52 249.685 12.57 249.815 ;
		RECT	13.98 249.685 14.03 249.815 ;
		RECT	14.33 402.555 14.38 402.685 ;
		RECT	6.22 403.015 6.27 403.145 ;
		RECT	7.5 403.015 7.55 403.145 ;
		RECT	9.04 403.015 9.09 403.145 ;
		RECT	9.315 403.015 9.365 403.145 ;
		RECT	9.72 403.015 9.77 403.145 ;
		RECT	11.025 403.015 11.075 403.145 ;
		RECT	12.79 403.015 12.84 403.145 ;
		RECT	14.33 404.975 14.38 405.105 ;
		RECT	5.675 405.205 5.725 405.335 ;
		RECT	6.065 405.205 6.115 405.335 ;
		RECT	6.725 405.205 6.775 405.335 ;
		RECT	8.42 405.205 8.47 405.335 ;
		RECT	8.77 405.205 8.82 405.335 ;
		RECT	11.555 405.205 11.605 405.335 ;
		RECT	11.815 405.205 11.865 405.335 ;
		RECT	12.52 405.205 12.57 405.335 ;
		RECT	13.98 405.205 14.03 405.335 ;
		RECT	14.33 405.435 14.38 405.565 ;
		RECT	6.22 405.895 6.27 406.025 ;
		RECT	7.5 405.895 7.55 406.025 ;
		RECT	9.04 405.895 9.09 406.025 ;
		RECT	9.315 405.895 9.365 406.025 ;
		RECT	9.72 405.895 9.77 406.025 ;
		RECT	11.025 405.895 11.075 406.025 ;
		RECT	12.79 405.895 12.84 406.025 ;
		RECT	14.33 407.855 14.38 407.985 ;
		RECT	5.675 408.085 5.725 408.215 ;
		RECT	6.065 408.085 6.115 408.215 ;
		RECT	6.725 408.085 6.775 408.215 ;
		RECT	8.42 408.085 8.47 408.215 ;
		RECT	8.77 408.085 8.82 408.215 ;
		RECT	11.555 408.085 11.605 408.215 ;
		RECT	11.815 408.085 11.865 408.215 ;
		RECT	12.52 408.085 12.57 408.215 ;
		RECT	13.98 408.085 14.03 408.215 ;
		RECT	14.33 408.315 14.38 408.445 ;
		RECT	6.22 408.775 6.27 408.905 ;
		RECT	7.5 408.775 7.55 408.905 ;
		RECT	9.04 408.775 9.09 408.905 ;
		RECT	9.315 408.775 9.365 408.905 ;
		RECT	9.72 408.775 9.77 408.905 ;
		RECT	11.025 408.775 11.075 408.905 ;
		RECT	12.79 408.775 12.84 408.905 ;
		RECT	14.33 410.735 14.38 410.865 ;
		RECT	5.675 410.965 5.725 411.095 ;
		RECT	6.065 410.965 6.115 411.095 ;
		RECT	6.725 410.965 6.775 411.095 ;
		RECT	8.42 410.965 8.47 411.095 ;
		RECT	8.77 410.965 8.82 411.095 ;
		RECT	11.555 410.965 11.605 411.095 ;
		RECT	11.815 410.965 11.865 411.095 ;
		RECT	12.52 410.965 12.57 411.095 ;
		RECT	13.98 410.965 14.03 411.095 ;
		RECT	14.33 249.915 14.38 250.045 ;
		RECT	6.22 250.375 6.27 250.505 ;
		RECT	7.5 250.375 7.55 250.505 ;
		RECT	9.04 250.375 9.09 250.505 ;
		RECT	9.315 250.375 9.365 250.505 ;
		RECT	9.72 250.375 9.77 250.505 ;
		RECT	11.025 250.375 11.075 250.505 ;
		RECT	12.79 250.375 12.84 250.505 ;
		RECT	14.33 252.335 14.38 252.465 ;
		RECT	5.675 252.565 5.725 252.695 ;
		RECT	6.065 252.565 6.115 252.695 ;
		RECT	6.725 252.565 6.775 252.695 ;
		RECT	8.42 252.565 8.47 252.695 ;
		RECT	8.77 252.565 8.82 252.695 ;
		RECT	11.555 252.565 11.605 252.695 ;
		RECT	11.815 252.565 11.865 252.695 ;
		RECT	12.52 252.565 12.57 252.695 ;
		RECT	13.98 252.565 14.03 252.695 ;
		RECT	14.33 252.795 14.38 252.925 ;
		RECT	6.22 253.255 6.27 253.385 ;
		RECT	7.5 253.255 7.55 253.385 ;
		RECT	9.04 253.255 9.09 253.385 ;
		RECT	9.315 253.255 9.365 253.385 ;
		RECT	9.72 253.255 9.77 253.385 ;
		RECT	11.025 253.255 11.075 253.385 ;
		RECT	12.79 253.255 12.84 253.385 ;
		RECT	14.33 255.215 14.38 255.345 ;
		RECT	5.675 255.445 5.725 255.575 ;
		RECT	6.065 255.445 6.115 255.575 ;
		RECT	6.725 255.445 6.775 255.575 ;
		RECT	8.42 255.445 8.47 255.575 ;
		RECT	8.77 255.445 8.82 255.575 ;
		RECT	11.555 255.445 11.605 255.575 ;
		RECT	11.815 255.445 11.865 255.575 ;
		RECT	12.52 255.445 12.57 255.575 ;
		RECT	13.98 255.445 14.03 255.575 ;
		RECT	14.33 255.675 14.38 255.805 ;
		RECT	6.22 256.135 6.27 256.265 ;
		RECT	7.5 256.135 7.55 256.265 ;
		RECT	9.04 256.135 9.09 256.265 ;
		RECT	9.315 256.135 9.365 256.265 ;
		RECT	9.72 256.135 9.77 256.265 ;
		RECT	11.025 256.135 11.075 256.265 ;
		RECT	12.79 256.135 12.84 256.265 ;
		RECT	14.33 258.095 14.38 258.225 ;
		RECT	5.675 258.325 5.725 258.455 ;
		RECT	6.065 258.325 6.115 258.455 ;
		RECT	6.725 258.325 6.775 258.455 ;
		RECT	8.42 258.325 8.47 258.455 ;
		RECT	8.77 258.325 8.82 258.455 ;
		RECT	11.555 258.325 11.605 258.455 ;
		RECT	11.815 258.325 11.865 258.455 ;
		RECT	12.52 258.325 12.57 258.455 ;
		RECT	13.98 258.325 14.03 258.455 ;
		RECT	14.33 411.195 14.38 411.325 ;
		RECT	6.22 411.655 6.27 411.785 ;
		RECT	7.5 411.655 7.55 411.785 ;
		RECT	9.04 411.655 9.09 411.785 ;
		RECT	9.315 411.655 9.365 411.785 ;
		RECT	9.72 411.655 9.77 411.785 ;
		RECT	11.025 411.655 11.075 411.785 ;
		RECT	12.79 411.655 12.84 411.785 ;
		RECT	14.33 413.615 14.38 413.745 ;
		RECT	5.675 413.845 5.725 413.975 ;
		RECT	6.065 413.845 6.115 413.975 ;
		RECT	6.725 413.845 6.775 413.975 ;
		RECT	8.42 413.845 8.47 413.975 ;
		RECT	8.77 413.845 8.82 413.975 ;
		RECT	11.555 413.845 11.605 413.975 ;
		RECT	11.815 413.845 11.865 413.975 ;
		RECT	12.52 413.845 12.57 413.975 ;
		RECT	13.98 413.845 14.03 413.975 ;
		RECT	14.33 229.755 14.38 229.885 ;
		RECT	6.22 230.215 6.27 230.345 ;
		RECT	7.5 230.215 7.55 230.345 ;
		RECT	9.04 230.215 9.09 230.345 ;
		RECT	9.315 230.215 9.365 230.345 ;
		RECT	9.72 230.215 9.77 230.345 ;
		RECT	11.025 230.215 11.075 230.345 ;
		RECT	12.79 230.215 12.84 230.345 ;
		RECT	14.33 232.175 14.38 232.305 ;
		RECT	5.675 232.405 5.725 232.535 ;
		RECT	6.065 232.405 6.115 232.535 ;
		RECT	6.725 232.405 6.775 232.535 ;
		RECT	8.42 232.405 8.47 232.535 ;
		RECT	8.77 232.405 8.82 232.535 ;
		RECT	11.555 232.405 11.605 232.535 ;
		RECT	11.815 232.405 11.865 232.535 ;
		RECT	12.52 232.405 12.57 232.535 ;
		RECT	13.98 232.405 14.03 232.535 ;
		RECT	13.98 414.535 14.03 414.665 ;
		RECT	3.06 414.075 3.11 414.205 ;
		RECT	1.57 414.535 1.62 414.665 ;
		RECT	2.485 414.535 2.665 414.665 ;
		RECT	3.84 414.535 3.89 414.665 ;
		RECT	7.19 414.535 7.24 414.665 ;
		RECT	14.14 414.535 14.19 414.665 ;
		RECT	13.8 414.305 13.85 414.435 ;
		RECT	8.56 414.075 8.61 414.205 ;
		RECT	10.27 414.075 10.32 414.205 ;
		RECT	0.435 414.075 0.485 414.205 ;
		RECT	0.62 414.535 0.67 414.665 ;
		RECT	3.65 414.535 3.7 414.665 ;
		RECT	2.18 414.075 2.23 414.205 ;
		RECT	0.9 235.285 0.95 235.415 ;
		RECT	0.9 261.205 0.95 261.335 ;
		RECT	0.9 264.085 0.95 264.215 ;
		RECT	0.9 266.965 0.95 267.095 ;
		RECT	0.9 269.845 0.95 269.975 ;
		RECT	0.9 272.725 0.95 272.855 ;
		RECT	0.9 275.605 0.95 275.735 ;
		RECT	0.9 278.485 0.95 278.615 ;
		RECT	0.9 281.365 0.95 281.495 ;
		RECT	0.9 284.245 0.95 284.375 ;
		RECT	0.9 287.125 0.95 287.255 ;
		RECT	0.9 238.165 0.95 238.295 ;
		RECT	0.9 290.005 0.95 290.135 ;
		RECT	0.9 292.885 0.95 293.015 ;
		RECT	0.9 295.765 0.95 295.895 ;
		RECT	0.9 298.645 0.95 298.775 ;
		RECT	0.9 301.525 0.95 301.655 ;
		RECT	0.9 304.405 0.95 304.535 ;
		RECT	0.9 307.285 0.95 307.415 ;
		RECT	0.9 310.165 0.95 310.295 ;
		RECT	0.9 313.045 0.95 313.175 ;
		RECT	0.9 315.925 0.95 316.055 ;
		RECT	0.9 241.045 0.95 241.175 ;
		RECT	0.9 318.805 0.95 318.935 ;
		RECT	0.9 321.685 0.95 321.815 ;
		RECT	0.9 324.565 0.95 324.695 ;
		RECT	0.9 327.445 0.95 327.575 ;
		RECT	0.9 330.325 0.95 330.455 ;
		RECT	0.9 333.205 0.95 333.335 ;
		RECT	0.9 336.085 0.95 336.215 ;
		RECT	0.9 338.965 0.95 339.095 ;
		RECT	0.9 341.845 0.95 341.975 ;
		RECT	0.9 344.725 0.95 344.855 ;
		RECT	0.9 243.925 0.95 244.055 ;
		RECT	0.9 347.605 0.95 347.735 ;
		RECT	0.9 350.485 0.95 350.615 ;
		RECT	0.9 353.365 0.95 353.495 ;
		RECT	0.9 356.245 0.95 356.375 ;
		RECT	0.9 359.125 0.95 359.255 ;
		RECT	0.9 362.005 0.95 362.135 ;
		RECT	0.9 364.885 0.95 365.015 ;
		RECT	0.9 367.765 0.95 367.895 ;
		RECT	0.9 370.645 0.95 370.775 ;
		RECT	0.9 373.525 0.95 373.655 ;
		RECT	0.9 246.805 0.95 246.935 ;
		RECT	0.9 376.405 0.95 376.535 ;
		RECT	0.9 379.285 0.95 379.415 ;
		RECT	0.9 382.165 0.95 382.295 ;
		RECT	0.9 385.045 0.95 385.175 ;
		RECT	0.9 387.925 0.95 388.055 ;
		RECT	0.9 390.805 0.95 390.935 ;
		RECT	0.9 393.685 0.95 393.815 ;
		RECT	0.9 396.565 0.95 396.695 ;
		RECT	0.9 399.445 0.95 399.575 ;
		RECT	0.9 402.325 0.95 402.455 ;
		RECT	0.9 249.685 0.95 249.815 ;
		RECT	0.9 405.205 0.95 405.335 ;
		RECT	0.9 408.085 0.95 408.215 ;
		RECT	0.9 410.965 0.95 411.095 ;
		RECT	0.9 252.565 0.95 252.695 ;
		RECT	0.9 255.445 0.95 255.575 ;
		RECT	0.9 258.325 0.95 258.455 ;
		RECT	0.9 413.845 0.95 413.975 ;
		RECT	0.9 232.405 0.95 232.535 ;
		RECT	2.18 229.755 2.23 229.885 ;
		RECT	2.18 232.175 2.23 232.305 ;
		RECT	2.18 258.555 2.23 258.685 ;
		RECT	2.18 260.975 2.23 261.105 ;
		RECT	2.18 261.435 2.23 261.565 ;
		RECT	2.18 263.855 2.23 263.985 ;
		RECT	2.18 264.315 2.23 264.445 ;
		RECT	2.18 266.735 2.23 266.865 ;
		RECT	2.18 267.195 2.23 267.325 ;
		RECT	2.18 269.615 2.23 269.745 ;
		RECT	2.18 270.075 2.23 270.205 ;
		RECT	2.18 272.495 2.23 272.625 ;
		RECT	2.18 272.955 2.23 273.085 ;
		RECT	2.18 275.375 2.23 275.505 ;
		RECT	2.18 275.835 2.23 275.965 ;
		RECT	2.18 278.255 2.23 278.385 ;
		RECT	2.18 278.715 2.23 278.845 ;
		RECT	2.18 281.135 2.23 281.265 ;
		RECT	2.18 281.595 2.23 281.725 ;
		RECT	2.18 284.015 2.23 284.145 ;
		RECT	2.18 284.475 2.23 284.605 ;
		RECT	2.18 286.895 2.23 287.025 ;
		RECT	2.18 232.635 2.23 232.765 ;
		RECT	2.18 235.055 2.23 235.185 ;
		RECT	2.18 287.355 2.23 287.485 ;
		RECT	2.18 289.775 2.23 289.905 ;
		RECT	2.18 290.235 2.23 290.365 ;
		RECT	2.18 292.655 2.23 292.785 ;
		RECT	2.18 293.115 2.23 293.245 ;
		RECT	2.18 295.535 2.23 295.665 ;
		RECT	2.18 295.995 2.23 296.125 ;
		RECT	2.18 298.415 2.23 298.545 ;
		RECT	2.18 298.875 2.23 299.005 ;
		RECT	2.18 301.295 2.23 301.425 ;
		RECT	2.18 301.755 2.23 301.885 ;
		RECT	2.18 304.175 2.23 304.305 ;
		RECT	2.18 304.635 2.23 304.765 ;
		RECT	2.18 307.055 2.23 307.185 ;
		RECT	2.18 307.515 2.23 307.645 ;
		RECT	2.18 309.935 2.23 310.065 ;
		RECT	2.18 310.395 2.23 310.525 ;
		RECT	2.18 312.815 2.23 312.945 ;
		RECT	2.18 313.275 2.23 313.405 ;
		RECT	2.18 315.695 2.23 315.825 ;
		RECT	2.18 235.515 2.23 235.645 ;
		RECT	2.18 237.935 2.23 238.065 ;
		RECT	2.18 316.155 2.23 316.285 ;
		RECT	2.18 318.575 2.23 318.705 ;
		RECT	2.18 319.035 2.23 319.165 ;
		RECT	2.18 321.455 2.23 321.585 ;
		RECT	2.18 321.915 2.23 322.045 ;
		RECT	2.18 324.335 2.23 324.465 ;
		RECT	2.18 324.795 2.23 324.925 ;
		RECT	2.18 327.215 2.23 327.345 ;
		RECT	2.18 327.675 2.23 327.805 ;
		RECT	2.18 330.095 2.23 330.225 ;
		RECT	2.18 330.555 2.23 330.685 ;
		RECT	2.18 332.975 2.23 333.105 ;
		RECT	2.18 333.435 2.23 333.565 ;
		RECT	2.18 335.855 2.23 335.985 ;
		RECT	2.18 336.315 2.23 336.445 ;
		RECT	2.18 338.735 2.23 338.865 ;
		RECT	2.18 339.195 2.23 339.325 ;
		RECT	2.18 341.615 2.23 341.745 ;
		RECT	2.18 342.075 2.23 342.205 ;
		RECT	2.18 344.495 2.23 344.625 ;
		RECT	2.18 238.395 2.23 238.525 ;
		RECT	2.18 240.815 2.23 240.945 ;
		RECT	2.18 344.955 2.23 345.085 ;
		RECT	2.18 347.375 2.23 347.505 ;
		RECT	2.18 347.835 2.23 347.965 ;
		RECT	2.18 350.255 2.23 350.385 ;
		RECT	2.18 350.715 2.23 350.845 ;
		RECT	2.18 353.135 2.23 353.265 ;
		RECT	2.18 353.595 2.23 353.725 ;
		RECT	2.18 356.015 2.23 356.145 ;
		RECT	2.18 356.475 2.23 356.605 ;
		RECT	2.18 358.895 2.23 359.025 ;
		RECT	2.18 359.355 2.23 359.485 ;
		RECT	2.18 361.775 2.23 361.905 ;
		RECT	2.18 362.235 2.23 362.365 ;
		RECT	2.18 364.655 2.23 364.785 ;
		RECT	2.18 365.115 2.23 365.245 ;
		RECT	2.18 367.535 2.23 367.665 ;
		RECT	2.18 367.995 2.23 368.125 ;
		RECT	2.18 370.415 2.23 370.545 ;
		RECT	2.18 370.875 2.23 371.005 ;
		RECT	2.18 373.295 2.23 373.425 ;
		RECT	2.18 241.275 2.23 241.405 ;
		RECT	2.18 243.695 2.23 243.825 ;
		RECT	2.18 373.755 2.23 373.885 ;
		RECT	2.18 376.175 2.23 376.305 ;
		RECT	2.18 376.635 2.23 376.765 ;
		RECT	2.18 379.055 2.23 379.185 ;
		RECT	2.18 379.515 2.23 379.645 ;
		RECT	2.18 381.935 2.23 382.065 ;
		RECT	2.18 382.395 2.23 382.525 ;
		RECT	2.18 384.815 2.23 384.945 ;
		RECT	2.18 385.275 2.23 385.405 ;
		RECT	2.18 387.695 2.23 387.825 ;
		RECT	2.18 388.155 2.23 388.285 ;
		RECT	2.18 390.575 2.23 390.705 ;
		RECT	2.18 391.035 2.23 391.165 ;
		RECT	2.18 393.455 2.23 393.585 ;
		RECT	2.18 393.915 2.23 394.045 ;
		RECT	2.18 396.335 2.23 396.465 ;
		RECT	2.18 396.795 2.23 396.925 ;
		RECT	2.18 399.215 2.23 399.345 ;
		RECT	2.18 399.675 2.23 399.805 ;
		RECT	2.18 402.095 2.23 402.225 ;
		RECT	2.18 244.155 2.23 244.285 ;
		RECT	2.18 246.575 2.23 246.705 ;
		RECT	2.18 402.555 2.23 402.685 ;
		RECT	2.18 404.975 2.23 405.105 ;
		RECT	2.18 405.435 2.23 405.565 ;
		RECT	2.18 407.855 2.23 407.985 ;
		RECT	2.18 408.315 2.23 408.445 ;
		RECT	2.18 410.735 2.23 410.865 ;
		RECT	2.18 411.195 2.23 411.325 ;
		RECT	2.18 413.615 2.23 413.745 ;
		RECT	2.18 247.035 2.23 247.165 ;
		RECT	2.18 249.455 2.23 249.585 ;
		RECT	2.18 249.915 2.23 250.045 ;
		RECT	2.18 252.335 2.23 252.465 ;
		RECT	2.18 252.795 2.23 252.925 ;
		RECT	2.18 255.215 2.23 255.345 ;
		RECT	2.18 255.675 2.23 255.805 ;
		RECT	2.18 258.095 2.23 258.225 ;
		RECT	1.38 229.755 1.43 229.885 ;
		RECT	4.51 229.755 4.56 229.885 ;
		RECT	3.06 230.215 3.11 230.345 ;
		RECT	1.405 232.175 1.455 232.305 ;
		RECT	4.51 232.175 4.56 232.305 ;
		RECT	1.38 258.555 1.43 258.685 ;
		RECT	4.51 258.555 4.56 258.685 ;
		RECT	3.06 259.015 3.11 259.145 ;
		RECT	1.405 260.975 1.455 261.105 ;
		RECT	4.51 260.975 4.56 261.105 ;
		RECT	1.38 261.435 1.43 261.565 ;
		RECT	4.51 261.435 4.56 261.565 ;
		RECT	3.06 261.895 3.11 262.025 ;
		RECT	1.405 263.855 1.455 263.985 ;
		RECT	4.51 263.855 4.56 263.985 ;
		RECT	1.38 264.315 1.43 264.445 ;
		RECT	4.51 264.315 4.56 264.445 ;
		RECT	3.06 264.775 3.11 264.905 ;
		RECT	1.405 266.735 1.455 266.865 ;
		RECT	4.51 266.735 4.56 266.865 ;
		RECT	1.38 267.195 1.43 267.325 ;
		RECT	4.51 267.195 4.56 267.325 ;
		RECT	3.06 267.655 3.11 267.785 ;
		RECT	1.405 269.615 1.455 269.745 ;
		RECT	4.51 269.615 4.56 269.745 ;
		RECT	1.38 270.075 1.43 270.205 ;
		RECT	4.51 270.075 4.56 270.205 ;
		RECT	3.06 270.535 3.11 270.665 ;
		RECT	1.405 272.495 1.455 272.625 ;
		RECT	4.51 272.495 4.56 272.625 ;
		RECT	1.38 272.955 1.43 273.085 ;
		RECT	4.51 272.955 4.56 273.085 ;
		RECT	3.06 273.415 3.11 273.545 ;
		RECT	1.405 275.375 1.455 275.505 ;
		RECT	4.51 275.375 4.56 275.505 ;
		RECT	1.38 275.835 1.43 275.965 ;
		RECT	4.51 275.835 4.56 275.965 ;
		RECT	3.06 276.295 3.11 276.425 ;
		RECT	1.405 278.255 1.455 278.385 ;
		RECT	4.51 278.255 4.56 278.385 ;
		RECT	1.38 278.715 1.43 278.845 ;
		RECT	4.51 278.715 4.56 278.845 ;
		RECT	3.06 279.175 3.11 279.305 ;
		RECT	1.405 281.135 1.455 281.265 ;
		RECT	4.51 281.135 4.56 281.265 ;
		RECT	1.38 281.595 1.43 281.725 ;
		RECT	4.51 281.595 4.56 281.725 ;
		RECT	3.06 282.055 3.11 282.185 ;
		RECT	1.405 284.015 1.455 284.145 ;
		RECT	4.51 284.015 4.56 284.145 ;
		RECT	1.38 284.475 1.43 284.605 ;
		RECT	4.51 284.475 4.56 284.605 ;
		RECT	3.06 284.935 3.11 285.065 ;
		RECT	1.405 286.895 1.455 287.025 ;
		RECT	4.51 286.895 4.56 287.025 ;
		RECT	1.38 232.635 1.43 232.765 ;
		RECT	4.51 232.635 4.56 232.765 ;
		RECT	3.06 233.095 3.11 233.225 ;
		RECT	1.405 235.055 1.455 235.185 ;
		RECT	4.51 235.055 4.56 235.185 ;
		RECT	1.38 287.355 1.43 287.485 ;
		RECT	4.51 287.355 4.56 287.485 ;
		RECT	3.06 287.815 3.11 287.945 ;
		RECT	1.405 289.775 1.455 289.905 ;
		RECT	4.51 289.775 4.56 289.905 ;
		RECT	1.38 290.235 1.43 290.365 ;
		RECT	4.51 290.235 4.56 290.365 ;
		RECT	3.06 290.695 3.11 290.825 ;
		RECT	1.405 292.655 1.455 292.785 ;
		RECT	4.51 292.655 4.56 292.785 ;
		RECT	1.38 293.115 1.43 293.245 ;
		RECT	4.51 293.115 4.56 293.245 ;
		RECT	3.06 293.575 3.11 293.705 ;
		RECT	1.405 295.535 1.455 295.665 ;
		RECT	4.51 295.535 4.56 295.665 ;
		RECT	1.38 295.995 1.43 296.125 ;
		RECT	4.51 295.995 4.56 296.125 ;
		RECT	3.06 296.455 3.11 296.585 ;
		RECT	1.405 298.415 1.455 298.545 ;
		RECT	4.51 298.415 4.56 298.545 ;
		RECT	1.38 298.875 1.43 299.005 ;
		RECT	4.51 298.875 4.56 299.005 ;
		RECT	3.06 299.335 3.11 299.465 ;
		RECT	1.405 301.295 1.455 301.425 ;
		RECT	4.51 301.295 4.56 301.425 ;
		RECT	1.38 301.755 1.43 301.885 ;
		RECT	4.51 301.755 4.56 301.885 ;
		RECT	3.06 302.215 3.11 302.345 ;
		RECT	1.405 304.175 1.455 304.305 ;
		RECT	4.51 304.175 4.56 304.305 ;
		RECT	1.38 304.635 1.43 304.765 ;
		RECT	4.51 304.635 4.56 304.765 ;
		RECT	3.06 305.095 3.11 305.225 ;
		RECT	1.405 307.055 1.455 307.185 ;
		RECT	4.51 307.055 4.56 307.185 ;
		RECT	1.38 307.515 1.43 307.645 ;
		RECT	4.51 307.515 4.56 307.645 ;
		RECT	3.06 307.975 3.11 308.105 ;
		RECT	1.405 309.935 1.455 310.065 ;
		RECT	4.51 309.935 4.56 310.065 ;
		RECT	1.38 310.395 1.43 310.525 ;
		RECT	4.51 310.395 4.56 310.525 ;
		RECT	3.06 310.855 3.11 310.985 ;
		RECT	1.405 312.815 1.455 312.945 ;
		RECT	4.51 312.815 4.56 312.945 ;
		RECT	1.38 313.275 1.43 313.405 ;
		RECT	4.51 313.275 4.56 313.405 ;
		RECT	3.06 313.735 3.11 313.865 ;
		RECT	1.405 315.695 1.455 315.825 ;
		RECT	4.51 315.695 4.56 315.825 ;
		RECT	1.38 235.515 1.43 235.645 ;
		RECT	4.51 235.515 4.56 235.645 ;
		RECT	3.06 235.975 3.11 236.105 ;
		RECT	1.405 237.935 1.455 238.065 ;
		RECT	4.51 237.935 4.56 238.065 ;
		RECT	1.38 316.155 1.43 316.285 ;
		RECT	4.51 316.155 4.56 316.285 ;
		RECT	3.06 316.615 3.11 316.745 ;
		RECT	1.405 318.575 1.455 318.705 ;
		RECT	4.51 318.575 4.56 318.705 ;
		RECT	1.38 319.035 1.43 319.165 ;
		RECT	4.51 319.035 4.56 319.165 ;
		RECT	3.06 319.495 3.11 319.625 ;
		RECT	1.405 321.455 1.455 321.585 ;
		RECT	4.51 321.455 4.56 321.585 ;
		RECT	1.38 321.915 1.43 322.045 ;
		RECT	4.51 321.915 4.56 322.045 ;
		RECT	3.06 322.375 3.11 322.505 ;
		RECT	1.405 324.335 1.455 324.465 ;
		RECT	4.51 324.335 4.56 324.465 ;
		RECT	1.38 324.795 1.43 324.925 ;
		RECT	4.51 324.795 4.56 324.925 ;
		RECT	3.06 325.255 3.11 325.385 ;
		RECT	1.405 327.215 1.455 327.345 ;
		RECT	4.51 327.215 4.56 327.345 ;
		RECT	1.38 327.675 1.43 327.805 ;
		RECT	4.51 327.675 4.56 327.805 ;
		RECT	3.06 328.135 3.11 328.265 ;
		RECT	1.405 330.095 1.455 330.225 ;
		RECT	4.51 330.095 4.56 330.225 ;
		RECT	1.38 330.555 1.43 330.685 ;
		RECT	4.51 330.555 4.56 330.685 ;
		RECT	3.06 331.015 3.11 331.145 ;
		RECT	1.405 332.975 1.455 333.105 ;
		RECT	4.51 332.975 4.56 333.105 ;
		RECT	1.38 333.435 1.43 333.565 ;
		RECT	4.51 333.435 4.56 333.565 ;
		RECT	3.06 333.895 3.11 334.025 ;
		RECT	1.405 335.855 1.455 335.985 ;
		RECT	4.51 335.855 4.56 335.985 ;
		RECT	1.38 336.315 1.43 336.445 ;
		RECT	4.51 336.315 4.56 336.445 ;
		RECT	3.06 336.775 3.11 336.905 ;
		RECT	1.405 338.735 1.455 338.865 ;
		RECT	4.51 338.735 4.56 338.865 ;
		RECT	1.38 339.195 1.43 339.325 ;
		RECT	4.51 339.195 4.56 339.325 ;
		RECT	3.06 339.655 3.11 339.785 ;
		RECT	1.405 341.615 1.455 341.745 ;
		RECT	4.51 341.615 4.56 341.745 ;
		RECT	1.38 342.075 1.43 342.205 ;
		RECT	4.51 342.075 4.56 342.205 ;
		RECT	3.06 342.535 3.11 342.665 ;
		RECT	1.405 344.495 1.455 344.625 ;
		RECT	4.51 344.495 4.56 344.625 ;
		RECT	1.38 238.395 1.43 238.525 ;
		RECT	4.51 238.395 4.56 238.525 ;
		RECT	3.06 238.855 3.11 238.985 ;
		RECT	1.405 240.815 1.455 240.945 ;
		RECT	4.51 240.815 4.56 240.945 ;
		RECT	1.38 344.955 1.43 345.085 ;
		RECT	4.51 344.955 4.56 345.085 ;
		RECT	3.06 345.415 3.11 345.545 ;
		RECT	1.405 347.375 1.455 347.505 ;
		RECT	4.51 347.375 4.56 347.505 ;
		RECT	1.38 347.835 1.43 347.965 ;
		RECT	4.51 347.835 4.56 347.965 ;
		RECT	3.06 348.295 3.11 348.425 ;
		RECT	1.405 350.255 1.455 350.385 ;
		RECT	4.51 350.255 4.56 350.385 ;
		RECT	1.38 350.715 1.43 350.845 ;
		RECT	4.51 350.715 4.56 350.845 ;
		RECT	3.06 351.175 3.11 351.305 ;
		RECT	1.405 353.135 1.455 353.265 ;
		RECT	4.51 353.135 4.56 353.265 ;
		RECT	1.38 353.595 1.43 353.725 ;
		RECT	4.51 353.595 4.56 353.725 ;
		RECT	3.06 354.055 3.11 354.185 ;
		RECT	1.405 356.015 1.455 356.145 ;
		RECT	4.51 356.015 4.56 356.145 ;
		RECT	1.38 356.475 1.43 356.605 ;
		RECT	4.51 356.475 4.56 356.605 ;
		RECT	3.06 356.935 3.11 357.065 ;
		RECT	1.405 358.895 1.455 359.025 ;
		RECT	4.51 358.895 4.56 359.025 ;
		RECT	1.38 359.355 1.43 359.485 ;
		RECT	4.51 359.355 4.56 359.485 ;
		RECT	3.06 359.815 3.11 359.945 ;
		RECT	1.405 361.775 1.455 361.905 ;
		RECT	4.51 361.775 4.56 361.905 ;
		RECT	1.38 362.235 1.43 362.365 ;
		RECT	4.51 362.235 4.56 362.365 ;
		RECT	3.06 362.695 3.11 362.825 ;
		RECT	1.405 364.655 1.455 364.785 ;
		RECT	4.51 364.655 4.56 364.785 ;
		RECT	1.38 365.115 1.43 365.245 ;
		RECT	4.51 365.115 4.56 365.245 ;
		RECT	3.06 365.575 3.11 365.705 ;
		RECT	1.405 367.535 1.455 367.665 ;
		RECT	4.51 367.535 4.56 367.665 ;
		RECT	1.38 367.995 1.43 368.125 ;
		RECT	4.51 367.995 4.56 368.125 ;
		RECT	3.06 368.455 3.11 368.585 ;
		RECT	1.405 370.415 1.455 370.545 ;
		RECT	4.51 370.415 4.56 370.545 ;
		RECT	1.38 370.875 1.43 371.005 ;
		RECT	4.51 370.875 4.56 371.005 ;
		RECT	3.06 371.335 3.11 371.465 ;
		RECT	1.405 373.295 1.455 373.425 ;
		RECT	4.51 373.295 4.56 373.425 ;
		RECT	1.38 241.275 1.43 241.405 ;
		RECT	4.51 241.275 4.56 241.405 ;
		RECT	3.06 241.735 3.11 241.865 ;
		RECT	1.405 243.695 1.455 243.825 ;
		RECT	4.51 243.695 4.56 243.825 ;
		RECT	1.38 373.755 1.43 373.885 ;
		RECT	4.51 373.755 4.56 373.885 ;
		RECT	3.06 374.215 3.11 374.345 ;
		RECT	1.405 376.175 1.455 376.305 ;
		RECT	4.51 376.175 4.56 376.305 ;
		RECT	1.38 376.635 1.43 376.765 ;
		RECT	4.51 376.635 4.56 376.765 ;
		RECT	3.06 377.095 3.11 377.225 ;
		RECT	1.405 379.055 1.455 379.185 ;
		RECT	4.51 379.055 4.56 379.185 ;
		RECT	1.38 379.515 1.43 379.645 ;
		RECT	4.51 379.515 4.56 379.645 ;
		RECT	3.06 379.975 3.11 380.105 ;
		RECT	1.405 381.935 1.455 382.065 ;
		RECT	4.51 381.935 4.56 382.065 ;
		RECT	1.38 382.395 1.43 382.525 ;
		RECT	4.51 382.395 4.56 382.525 ;
		RECT	3.06 382.855 3.11 382.985 ;
		RECT	1.405 384.815 1.455 384.945 ;
		RECT	4.51 384.815 4.56 384.945 ;
		RECT	1.38 385.275 1.43 385.405 ;
		RECT	4.51 385.275 4.56 385.405 ;
		RECT	3.06 385.735 3.11 385.865 ;
		RECT	1.405 387.695 1.455 387.825 ;
		RECT	4.51 387.695 4.56 387.825 ;
		RECT	1.38 388.155 1.43 388.285 ;
		RECT	4.51 388.155 4.56 388.285 ;
		RECT	3.06 388.615 3.11 388.745 ;
		RECT	1.405 390.575 1.455 390.705 ;
		RECT	4.51 390.575 4.56 390.705 ;
		RECT	1.38 391.035 1.43 391.165 ;
		RECT	4.51 391.035 4.56 391.165 ;
		RECT	3.06 391.495 3.11 391.625 ;
		RECT	1.405 393.455 1.455 393.585 ;
		RECT	4.51 393.455 4.56 393.585 ;
		RECT	1.38 393.915 1.43 394.045 ;
		RECT	4.51 393.915 4.56 394.045 ;
		RECT	3.06 394.375 3.11 394.505 ;
		RECT	1.405 396.335 1.455 396.465 ;
		RECT	4.51 396.335 4.56 396.465 ;
		RECT	1.38 396.795 1.43 396.925 ;
		RECT	4.51 396.795 4.56 396.925 ;
		RECT	3.06 397.255 3.11 397.385 ;
		RECT	1.405 399.215 1.455 399.345 ;
		RECT	4.51 399.215 4.56 399.345 ;
		RECT	1.38 399.675 1.43 399.805 ;
		RECT	4.51 399.675 4.56 399.805 ;
		RECT	3.06 400.135 3.11 400.265 ;
		RECT	1.405 402.095 1.455 402.225 ;
		RECT	4.51 402.095 4.56 402.225 ;
		RECT	1.38 244.155 1.43 244.285 ;
		RECT	4.51 244.155 4.56 244.285 ;
		RECT	3.06 244.615 3.11 244.745 ;
		RECT	1.405 246.575 1.455 246.705 ;
		RECT	4.51 246.575 4.56 246.705 ;
		RECT	1.38 402.555 1.43 402.685 ;
		RECT	4.51 402.555 4.56 402.685 ;
		RECT	3.06 403.015 3.11 403.145 ;
		RECT	1.405 404.975 1.455 405.105 ;
		RECT	4.51 404.975 4.56 405.105 ;
		RECT	1.38 405.435 1.43 405.565 ;
		RECT	4.51 405.435 4.56 405.565 ;
		RECT	3.06 405.895 3.11 406.025 ;
		RECT	1.405 407.855 1.455 407.985 ;
		RECT	4.51 407.855 4.56 407.985 ;
		RECT	1.38 408.315 1.43 408.445 ;
		RECT	4.51 408.315 4.56 408.445 ;
		RECT	3.06 408.775 3.11 408.905 ;
		RECT	1.405 410.735 1.455 410.865 ;
		RECT	4.51 410.735 4.56 410.865 ;
		RECT	1.38 411.195 1.43 411.325 ;
		RECT	4.51 411.195 4.56 411.325 ;
		RECT	3.06 411.655 3.11 411.785 ;
		RECT	1.405 413.615 1.455 413.745 ;
		RECT	4.51 413.615 4.56 413.745 ;
		RECT	1.38 247.035 1.43 247.165 ;
		RECT	4.51 247.035 4.56 247.165 ;
		RECT	3.06 247.495 3.11 247.625 ;
		RECT	1.405 249.455 1.455 249.585 ;
		RECT	4.51 249.455 4.56 249.585 ;
		RECT	1.38 249.915 1.43 250.045 ;
		RECT	4.51 249.915 4.56 250.045 ;
		RECT	3.06 250.375 3.11 250.505 ;
		RECT	1.405 252.335 1.455 252.465 ;
		RECT	4.51 252.335 4.56 252.465 ;
		RECT	1.38 252.795 1.43 252.925 ;
		RECT	4.51 252.795 4.56 252.925 ;
		RECT	3.06 253.255 3.11 253.385 ;
		RECT	1.405 255.215 1.455 255.345 ;
		RECT	4.51 255.215 4.56 255.345 ;
		RECT	1.38 255.675 1.43 255.805 ;
		RECT	4.51 255.675 4.56 255.805 ;
		RECT	3.06 256.135 3.11 256.265 ;
		RECT	1.405 258.095 1.455 258.225 ;
		RECT	4.51 258.095 4.56 258.225 ;
		RECT	3.06 232.635 3.11 232.765 ;
		RECT	1.085 233.095 1.135 233.225 ;
		RECT	1.405 233.135 1.455 233.185 ;
		RECT	4.47 233.135 4.6 233.185 ;
		RECT	3.06 235.055 3.11 235.185 ;
		RECT	1.57 235.285 1.62 235.415 ;
		RECT	2.58 235.285 2.63 235.415 ;
		RECT	3.84 235.285 3.89 235.415 ;
		RECT	5.675 235.285 5.725 235.415 ;
		RECT	3.06 258.555 3.11 258.685 ;
		RECT	1.085 259.015 1.135 259.145 ;
		RECT	1.405 259.055 1.455 259.105 ;
		RECT	4.47 259.055 4.6 259.105 ;
		RECT	3.06 260.975 3.11 261.105 ;
		RECT	1.57 261.205 1.62 261.335 ;
		RECT	2.58 261.205 2.63 261.335 ;
		RECT	3.84 261.205 3.89 261.335 ;
		RECT	5.675 261.205 5.725 261.335 ;
		RECT	3.06 261.435 3.11 261.565 ;
		RECT	1.085 261.895 1.135 262.025 ;
		RECT	1.405 261.935 1.455 261.985 ;
		RECT	4.47 261.935 4.6 261.985 ;
		RECT	3.06 263.855 3.11 263.985 ;
		RECT	1.57 264.085 1.62 264.215 ;
		RECT	2.58 264.085 2.63 264.215 ;
		RECT	3.84 264.085 3.89 264.215 ;
		RECT	5.675 264.085 5.725 264.215 ;
		RECT	3.06 264.315 3.11 264.445 ;
		RECT	1.085 264.775 1.135 264.905 ;
		RECT	1.405 264.815 1.455 264.865 ;
		RECT	4.47 264.815 4.6 264.865 ;
		RECT	3.06 266.735 3.11 266.865 ;
		RECT	1.57 266.965 1.62 267.095 ;
		RECT	2.58 266.965 2.63 267.095 ;
		RECT	3.84 266.965 3.89 267.095 ;
		RECT	5.675 266.965 5.725 267.095 ;
		RECT	3.06 267.195 3.11 267.325 ;
		RECT	1.085 267.655 1.135 267.785 ;
		RECT	1.405 267.695 1.455 267.745 ;
		RECT	4.47 267.695 4.6 267.745 ;
		RECT	3.06 269.615 3.11 269.745 ;
		RECT	1.57 269.845 1.62 269.975 ;
		RECT	2.58 269.845 2.63 269.975 ;
		RECT	3.84 269.845 3.89 269.975 ;
		RECT	5.675 269.845 5.725 269.975 ;
		RECT	3.06 270.075 3.11 270.205 ;
		RECT	1.085 270.535 1.135 270.665 ;
		RECT	1.405 270.575 1.455 270.625 ;
		RECT	4.47 270.575 4.6 270.625 ;
		RECT	3.06 272.495 3.11 272.625 ;
		RECT	1.57 272.725 1.62 272.855 ;
		RECT	2.58 272.725 2.63 272.855 ;
		RECT	3.84 272.725 3.89 272.855 ;
		RECT	5.675 272.725 5.725 272.855 ;
		RECT	3.06 272.955 3.11 273.085 ;
		RECT	1.085 273.415 1.135 273.545 ;
		RECT	1.405 273.455 1.455 273.505 ;
		RECT	4.47 273.455 4.6 273.505 ;
		RECT	3.06 275.375 3.11 275.505 ;
		RECT	1.57 275.605 1.62 275.735 ;
		RECT	2.58 275.605 2.63 275.735 ;
		RECT	3.84 275.605 3.89 275.735 ;
		RECT	5.675 275.605 5.725 275.735 ;
		RECT	3.06 275.835 3.11 275.965 ;
		RECT	1.085 276.295 1.135 276.425 ;
		RECT	1.405 276.335 1.455 276.385 ;
		RECT	4.47 276.335 4.6 276.385 ;
		RECT	3.06 278.255 3.11 278.385 ;
		RECT	1.57 278.485 1.62 278.615 ;
		RECT	2.58 278.485 2.63 278.615 ;
		RECT	3.84 278.485 3.89 278.615 ;
		RECT	5.675 278.485 5.725 278.615 ;
		RECT	3.06 278.715 3.11 278.845 ;
		RECT	1.085 279.175 1.135 279.305 ;
		RECT	1.405 279.215 1.455 279.265 ;
		RECT	4.47 279.215 4.6 279.265 ;
		RECT	3.06 281.135 3.11 281.265 ;
		RECT	1.57 281.365 1.62 281.495 ;
		RECT	2.58 281.365 2.63 281.495 ;
		RECT	3.84 281.365 3.89 281.495 ;
		RECT	5.675 281.365 5.725 281.495 ;
		RECT	3.06 281.595 3.11 281.725 ;
		RECT	1.085 282.055 1.135 282.185 ;
		RECT	1.405 282.095 1.455 282.145 ;
		RECT	4.47 282.095 4.6 282.145 ;
		RECT	3.06 284.015 3.11 284.145 ;
		RECT	1.57 284.245 1.62 284.375 ;
		RECT	2.58 284.245 2.63 284.375 ;
		RECT	3.84 284.245 3.89 284.375 ;
		RECT	5.675 284.245 5.725 284.375 ;
		RECT	3.06 284.475 3.11 284.605 ;
		RECT	1.085 284.935 1.135 285.065 ;
		RECT	1.405 284.975 1.455 285.025 ;
		RECT	4.47 284.975 4.6 285.025 ;
		RECT	3.06 286.895 3.11 287.025 ;
		RECT	1.57 287.125 1.62 287.255 ;
		RECT	2.58 287.125 2.63 287.255 ;
		RECT	3.84 287.125 3.89 287.255 ;
		RECT	5.675 287.125 5.725 287.255 ;
		RECT	3.06 235.515 3.11 235.645 ;
		RECT	1.085 235.975 1.135 236.105 ;
		RECT	1.405 236.015 1.455 236.065 ;
		RECT	4.47 236.015 4.6 236.065 ;
		RECT	3.06 237.935 3.11 238.065 ;
		RECT	1.57 238.165 1.62 238.295 ;
		RECT	2.58 238.165 2.63 238.295 ;
		RECT	3.84 238.165 3.89 238.295 ;
		RECT	5.675 238.165 5.725 238.295 ;
		RECT	3.06 287.355 3.11 287.485 ;
		RECT	1.085 287.815 1.135 287.945 ;
		RECT	1.405 287.855 1.455 287.905 ;
		RECT	4.47 287.855 4.6 287.905 ;
		RECT	3.06 289.775 3.11 289.905 ;
		RECT	1.57 290.005 1.62 290.135 ;
		RECT	2.58 290.005 2.63 290.135 ;
		RECT	3.84 290.005 3.89 290.135 ;
		RECT	5.675 290.005 5.725 290.135 ;
		RECT	3.06 290.235 3.11 290.365 ;
		RECT	1.085 290.695 1.135 290.825 ;
		RECT	1.405 290.735 1.455 290.785 ;
		RECT	4.47 290.735 4.6 290.785 ;
		RECT	3.06 292.655 3.11 292.785 ;
		RECT	1.57 292.885 1.62 293.015 ;
		RECT	2.58 292.885 2.63 293.015 ;
		RECT	3.84 292.885 3.89 293.015 ;
		RECT	5.675 292.885 5.725 293.015 ;
		RECT	3.06 293.115 3.11 293.245 ;
		RECT	1.085 293.575 1.135 293.705 ;
		RECT	1.405 293.615 1.455 293.665 ;
		RECT	4.47 293.615 4.6 293.665 ;
		RECT	3.06 295.535 3.11 295.665 ;
		RECT	1.57 295.765 1.62 295.895 ;
		RECT	2.58 295.765 2.63 295.895 ;
		RECT	3.84 295.765 3.89 295.895 ;
		RECT	5.675 295.765 5.725 295.895 ;
		RECT	3.06 295.995 3.11 296.125 ;
		RECT	1.085 296.455 1.135 296.585 ;
		RECT	1.405 296.495 1.455 296.545 ;
		RECT	4.47 296.495 4.6 296.545 ;
		RECT	3.06 298.415 3.11 298.545 ;
		RECT	1.57 298.645 1.62 298.775 ;
		RECT	2.58 298.645 2.63 298.775 ;
		RECT	3.84 298.645 3.89 298.775 ;
		RECT	5.675 298.645 5.725 298.775 ;
		RECT	3.06 298.875 3.11 299.005 ;
		RECT	1.085 299.335 1.135 299.465 ;
		RECT	1.405 299.375 1.455 299.425 ;
		RECT	4.47 299.375 4.6 299.425 ;
		RECT	3.06 301.295 3.11 301.425 ;
		RECT	1.57 301.525 1.62 301.655 ;
		RECT	2.58 301.525 2.63 301.655 ;
		RECT	3.84 301.525 3.89 301.655 ;
		RECT	5.675 301.525 5.725 301.655 ;
		RECT	3.06 301.755 3.11 301.885 ;
		RECT	1.085 302.215 1.135 302.345 ;
		RECT	1.405 302.255 1.455 302.305 ;
		RECT	4.47 302.255 4.6 302.305 ;
		RECT	3.06 304.175 3.11 304.305 ;
		RECT	1.57 304.405 1.62 304.535 ;
		RECT	2.58 304.405 2.63 304.535 ;
		RECT	3.84 304.405 3.89 304.535 ;
		RECT	5.675 304.405 5.725 304.535 ;
		RECT	3.06 304.635 3.11 304.765 ;
		RECT	1.085 305.095 1.135 305.225 ;
		RECT	1.405 305.135 1.455 305.185 ;
		RECT	4.47 305.135 4.6 305.185 ;
		RECT	3.06 307.055 3.11 307.185 ;
		RECT	1.57 307.285 1.62 307.415 ;
		RECT	2.58 307.285 2.63 307.415 ;
		RECT	3.84 307.285 3.89 307.415 ;
		RECT	5.675 307.285 5.725 307.415 ;
		RECT	3.06 307.515 3.11 307.645 ;
		RECT	1.085 307.975 1.135 308.105 ;
		RECT	1.405 308.015 1.455 308.065 ;
		RECT	4.47 308.015 4.6 308.065 ;
		RECT	3.06 309.935 3.11 310.065 ;
		RECT	1.57 310.165 1.62 310.295 ;
		RECT	2.58 310.165 2.63 310.295 ;
		RECT	3.84 310.165 3.89 310.295 ;
		RECT	5.675 310.165 5.725 310.295 ;
		RECT	3.06 310.395 3.11 310.525 ;
		RECT	1.085 310.855 1.135 310.985 ;
		RECT	1.405 310.895 1.455 310.945 ;
		RECT	4.47 310.895 4.6 310.945 ;
		RECT	3.06 312.815 3.11 312.945 ;
		RECT	1.57 313.045 1.62 313.175 ;
		RECT	2.58 313.045 2.63 313.175 ;
		RECT	3.84 313.045 3.89 313.175 ;
		RECT	5.675 313.045 5.725 313.175 ;
		RECT	3.06 313.275 3.11 313.405 ;
		RECT	1.085 313.735 1.135 313.865 ;
		RECT	1.405 313.775 1.455 313.825 ;
		RECT	4.47 313.775 4.6 313.825 ;
		RECT	3.06 315.695 3.11 315.825 ;
		RECT	1.57 315.925 1.62 316.055 ;
		RECT	2.58 315.925 2.63 316.055 ;
		RECT	3.84 315.925 3.89 316.055 ;
		RECT	5.675 315.925 5.725 316.055 ;
		RECT	3.06 238.395 3.11 238.525 ;
		RECT	1.085 238.855 1.135 238.985 ;
		RECT	1.405 238.895 1.455 238.945 ;
		RECT	4.47 238.895 4.6 238.945 ;
		RECT	3.06 240.815 3.11 240.945 ;
		RECT	1.57 241.045 1.62 241.175 ;
		RECT	2.58 241.045 2.63 241.175 ;
		RECT	3.84 241.045 3.89 241.175 ;
		RECT	5.675 241.045 5.725 241.175 ;
		RECT	3.06 316.155 3.11 316.285 ;
		RECT	1.085 316.615 1.135 316.745 ;
		RECT	1.405 316.655 1.455 316.705 ;
		RECT	4.47 316.655 4.6 316.705 ;
		RECT	3.06 318.575 3.11 318.705 ;
		RECT	1.57 318.805 1.62 318.935 ;
		RECT	2.58 318.805 2.63 318.935 ;
		RECT	3.84 318.805 3.89 318.935 ;
		RECT	5.675 318.805 5.725 318.935 ;
		RECT	3.06 319.035 3.11 319.165 ;
		RECT	1.085 319.495 1.135 319.625 ;
		RECT	1.405 319.535 1.455 319.585 ;
		RECT	4.47 319.535 4.6 319.585 ;
		RECT	3.06 321.455 3.11 321.585 ;
		RECT	1.57 321.685 1.62 321.815 ;
		RECT	2.58 321.685 2.63 321.815 ;
		RECT	3.84 321.685 3.89 321.815 ;
		RECT	5.675 321.685 5.725 321.815 ;
		RECT	3.06 321.915 3.11 322.045 ;
		RECT	1.085 322.375 1.135 322.505 ;
		RECT	1.405 322.415 1.455 322.465 ;
		RECT	4.47 322.415 4.6 322.465 ;
		RECT	3.06 324.335 3.11 324.465 ;
		RECT	1.57 324.565 1.62 324.695 ;
		RECT	2.58 324.565 2.63 324.695 ;
		RECT	3.84 324.565 3.89 324.695 ;
		RECT	5.675 324.565 5.725 324.695 ;
		RECT	3.06 324.795 3.11 324.925 ;
		RECT	1.085 325.255 1.135 325.385 ;
		RECT	1.405 325.295 1.455 325.345 ;
		RECT	4.47 325.295 4.6 325.345 ;
		RECT	3.06 327.215 3.11 327.345 ;
		RECT	1.57 327.445 1.62 327.575 ;
		RECT	2.58 327.445 2.63 327.575 ;
		RECT	3.84 327.445 3.89 327.575 ;
		RECT	5.675 327.445 5.725 327.575 ;
		RECT	3.06 327.675 3.11 327.805 ;
		RECT	1.085 328.135 1.135 328.265 ;
		RECT	1.405 328.175 1.455 328.225 ;
		RECT	4.47 328.175 4.6 328.225 ;
		RECT	3.06 330.095 3.11 330.225 ;
		RECT	1.57 330.325 1.62 330.455 ;
		RECT	2.58 330.325 2.63 330.455 ;
		RECT	3.84 330.325 3.89 330.455 ;
		RECT	5.675 330.325 5.725 330.455 ;
		RECT	3.06 330.555 3.11 330.685 ;
		RECT	1.085 331.015 1.135 331.145 ;
		RECT	1.405 331.055 1.455 331.105 ;
		RECT	4.47 331.055 4.6 331.105 ;
		RECT	3.06 332.975 3.11 333.105 ;
		RECT	1.57 333.205 1.62 333.335 ;
		RECT	2.58 333.205 2.63 333.335 ;
		RECT	3.84 333.205 3.89 333.335 ;
		RECT	5.675 333.205 5.725 333.335 ;
		RECT	3.06 333.435 3.11 333.565 ;
		RECT	1.085 333.895 1.135 334.025 ;
		RECT	1.405 333.935 1.455 333.985 ;
		RECT	4.47 333.935 4.6 333.985 ;
		RECT	3.06 335.855 3.11 335.985 ;
		RECT	1.57 336.085 1.62 336.215 ;
		RECT	2.58 336.085 2.63 336.215 ;
		RECT	3.84 336.085 3.89 336.215 ;
		RECT	5.675 336.085 5.725 336.215 ;
		RECT	3.06 336.315 3.11 336.445 ;
		RECT	1.085 336.775 1.135 336.905 ;
		RECT	1.405 336.815 1.455 336.865 ;
		RECT	4.47 336.815 4.6 336.865 ;
		RECT	3.06 338.735 3.11 338.865 ;
		RECT	1.57 338.965 1.62 339.095 ;
		RECT	2.58 338.965 2.63 339.095 ;
		RECT	3.84 338.965 3.89 339.095 ;
		RECT	5.675 338.965 5.725 339.095 ;
		RECT	3.06 339.195 3.11 339.325 ;
		RECT	1.085 339.655 1.135 339.785 ;
		RECT	1.405 339.695 1.455 339.745 ;
		RECT	4.47 339.695 4.6 339.745 ;
		RECT	3.06 341.615 3.11 341.745 ;
		RECT	1.57 341.845 1.62 341.975 ;
		RECT	2.58 341.845 2.63 341.975 ;
		RECT	3.84 341.845 3.89 341.975 ;
		RECT	5.675 341.845 5.725 341.975 ;
		RECT	3.06 342.075 3.11 342.205 ;
		RECT	1.085 342.535 1.135 342.665 ;
		RECT	1.405 342.575 1.455 342.625 ;
		RECT	4.47 342.575 4.6 342.625 ;
		RECT	3.06 344.495 3.11 344.625 ;
		RECT	1.57 344.725 1.62 344.855 ;
		RECT	2.58 344.725 2.63 344.855 ;
		RECT	3.84 344.725 3.89 344.855 ;
		RECT	5.675 344.725 5.725 344.855 ;
		RECT	3.06 241.275 3.11 241.405 ;
		RECT	1.085 241.735 1.135 241.865 ;
		RECT	1.405 241.775 1.455 241.825 ;
		RECT	4.47 241.775 4.6 241.825 ;
		RECT	3.06 243.695 3.11 243.825 ;
		RECT	1.57 243.925 1.62 244.055 ;
		RECT	2.58 243.925 2.63 244.055 ;
		RECT	3.84 243.925 3.89 244.055 ;
		RECT	5.675 243.925 5.725 244.055 ;
		RECT	3.06 344.955 3.11 345.085 ;
		RECT	1.085 345.415 1.135 345.545 ;
		RECT	1.405 345.455 1.455 345.505 ;
		RECT	4.47 345.455 4.6 345.505 ;
		RECT	3.06 347.375 3.11 347.505 ;
		RECT	1.57 347.605 1.62 347.735 ;
		RECT	2.58 347.605 2.63 347.735 ;
		RECT	3.84 347.605 3.89 347.735 ;
		RECT	5.675 347.605 5.725 347.735 ;
		RECT	3.06 347.835 3.11 347.965 ;
		RECT	1.085 348.295 1.135 348.425 ;
		RECT	1.405 348.335 1.455 348.385 ;
		RECT	4.47 348.335 4.6 348.385 ;
		RECT	3.06 350.255 3.11 350.385 ;
		RECT	1.57 350.485 1.62 350.615 ;
		RECT	2.58 350.485 2.63 350.615 ;
		RECT	3.84 350.485 3.89 350.615 ;
		RECT	5.675 350.485 5.725 350.615 ;
		RECT	3.06 350.715 3.11 350.845 ;
		RECT	1.085 351.175 1.135 351.305 ;
		RECT	1.405 351.215 1.455 351.265 ;
		RECT	4.47 351.215 4.6 351.265 ;
		RECT	3.06 353.135 3.11 353.265 ;
		RECT	1.57 353.365 1.62 353.495 ;
		RECT	2.58 353.365 2.63 353.495 ;
		RECT	3.84 353.365 3.89 353.495 ;
		RECT	5.675 353.365 5.725 353.495 ;
		RECT	3.06 353.595 3.11 353.725 ;
		RECT	1.085 354.055 1.135 354.185 ;
		RECT	1.405 354.095 1.455 354.145 ;
		RECT	4.47 354.095 4.6 354.145 ;
		RECT	3.06 356.015 3.11 356.145 ;
		RECT	1.57 356.245 1.62 356.375 ;
		RECT	2.58 356.245 2.63 356.375 ;
		RECT	3.84 356.245 3.89 356.375 ;
		RECT	5.675 356.245 5.725 356.375 ;
		RECT	3.06 356.475 3.11 356.605 ;
		RECT	1.085 356.935 1.135 357.065 ;
		RECT	1.405 356.975 1.455 357.025 ;
		RECT	4.47 356.975 4.6 357.025 ;
		RECT	3.06 358.895 3.11 359.025 ;
		RECT	1.57 359.125 1.62 359.255 ;
		RECT	2.58 359.125 2.63 359.255 ;
		RECT	3.84 359.125 3.89 359.255 ;
		RECT	5.675 359.125 5.725 359.255 ;
		RECT	3.06 359.355 3.11 359.485 ;
		RECT	1.085 359.815 1.135 359.945 ;
		RECT	1.405 359.855 1.455 359.905 ;
		RECT	4.47 359.855 4.6 359.905 ;
		RECT	3.06 361.775 3.11 361.905 ;
		RECT	1.57 362.005 1.62 362.135 ;
		RECT	2.58 362.005 2.63 362.135 ;
		RECT	3.84 362.005 3.89 362.135 ;
		RECT	5.675 362.005 5.725 362.135 ;
		RECT	3.06 362.235 3.11 362.365 ;
		RECT	1.085 362.695 1.135 362.825 ;
		RECT	1.405 362.735 1.455 362.785 ;
		RECT	4.47 362.735 4.6 362.785 ;
		RECT	3.06 364.655 3.11 364.785 ;
		RECT	1.57 364.885 1.62 365.015 ;
		RECT	2.58 364.885 2.63 365.015 ;
		RECT	3.84 364.885 3.89 365.015 ;
		RECT	5.675 364.885 5.725 365.015 ;
		RECT	3.06 365.115 3.11 365.245 ;
		RECT	1.085 365.575 1.135 365.705 ;
		RECT	1.405 365.615 1.455 365.665 ;
		RECT	4.47 365.615 4.6 365.665 ;
		RECT	3.06 367.535 3.11 367.665 ;
		RECT	1.57 367.765 1.62 367.895 ;
		RECT	2.58 367.765 2.63 367.895 ;
		RECT	3.84 367.765 3.89 367.895 ;
		RECT	5.675 367.765 5.725 367.895 ;
		RECT	3.06 367.995 3.11 368.125 ;
		RECT	1.085 368.455 1.135 368.585 ;
		RECT	1.405 368.495 1.455 368.545 ;
		RECT	4.47 368.495 4.6 368.545 ;
		RECT	3.06 370.415 3.11 370.545 ;
		RECT	1.57 370.645 1.62 370.775 ;
		RECT	2.58 370.645 2.63 370.775 ;
		RECT	3.84 370.645 3.89 370.775 ;
		RECT	5.675 370.645 5.725 370.775 ;
		RECT	3.06 370.875 3.11 371.005 ;
		RECT	1.085 371.335 1.135 371.465 ;
		RECT	1.405 371.375 1.455 371.425 ;
		RECT	4.47 371.375 4.6 371.425 ;
		RECT	3.06 373.295 3.11 373.425 ;
		RECT	1.57 373.525 1.62 373.655 ;
		RECT	2.58 373.525 2.63 373.655 ;
		RECT	3.84 373.525 3.89 373.655 ;
		RECT	5.675 373.525 5.725 373.655 ;
		RECT	3.06 244.155 3.11 244.285 ;
		RECT	1.085 244.615 1.135 244.745 ;
		RECT	1.405 244.655 1.455 244.705 ;
		RECT	4.47 244.655 4.6 244.705 ;
		RECT	3.06 246.575 3.11 246.705 ;
		RECT	1.57 246.805 1.62 246.935 ;
		RECT	2.58 246.805 2.63 246.935 ;
		RECT	3.84 246.805 3.89 246.935 ;
		RECT	5.675 246.805 5.725 246.935 ;
		RECT	3.06 373.755 3.11 373.885 ;
		RECT	1.085 374.215 1.135 374.345 ;
		RECT	1.405 374.255 1.455 374.305 ;
		RECT	4.47 374.255 4.6 374.305 ;
		RECT	3.06 376.175 3.11 376.305 ;
		RECT	1.57 376.405 1.62 376.535 ;
		RECT	2.58 376.405 2.63 376.535 ;
		RECT	3.84 376.405 3.89 376.535 ;
		RECT	5.675 376.405 5.725 376.535 ;
		RECT	3.06 376.635 3.11 376.765 ;
		RECT	1.085 377.095 1.135 377.225 ;
		RECT	1.405 377.135 1.455 377.185 ;
		RECT	4.47 377.135 4.6 377.185 ;
		RECT	3.06 379.055 3.11 379.185 ;
		RECT	1.57 379.285 1.62 379.415 ;
		RECT	2.58 379.285 2.63 379.415 ;
		RECT	3.84 379.285 3.89 379.415 ;
		RECT	5.675 379.285 5.725 379.415 ;
		RECT	3.06 379.515 3.11 379.645 ;
		RECT	1.085 379.975 1.135 380.105 ;
		RECT	1.405 380.015 1.455 380.065 ;
		RECT	4.47 380.015 4.6 380.065 ;
		RECT	3.06 381.935 3.11 382.065 ;
		RECT	1.57 382.165 1.62 382.295 ;
		RECT	2.58 382.165 2.63 382.295 ;
		RECT	3.84 382.165 3.89 382.295 ;
		RECT	5.675 382.165 5.725 382.295 ;
		RECT	3.06 382.395 3.11 382.525 ;
		RECT	1.085 382.855 1.135 382.985 ;
		RECT	1.405 382.895 1.455 382.945 ;
		RECT	4.47 382.895 4.6 382.945 ;
		RECT	3.06 384.815 3.11 384.945 ;
		RECT	1.57 385.045 1.62 385.175 ;
		RECT	2.58 385.045 2.63 385.175 ;
		RECT	3.84 385.045 3.89 385.175 ;
		RECT	5.675 385.045 5.725 385.175 ;
		RECT	3.06 385.275 3.11 385.405 ;
		RECT	1.085 385.735 1.135 385.865 ;
		RECT	1.405 385.775 1.455 385.825 ;
		RECT	4.47 385.775 4.6 385.825 ;
		RECT	3.06 387.695 3.11 387.825 ;
		RECT	1.57 387.925 1.62 388.055 ;
		RECT	2.58 387.925 2.63 388.055 ;
		RECT	3.84 387.925 3.89 388.055 ;
		RECT	5.675 387.925 5.725 388.055 ;
		RECT	3.06 388.155 3.11 388.285 ;
		RECT	1.085 388.615 1.135 388.745 ;
		RECT	1.405 388.655 1.455 388.705 ;
		RECT	4.47 388.655 4.6 388.705 ;
		RECT	3.06 390.575 3.11 390.705 ;
		RECT	1.57 390.805 1.62 390.935 ;
		RECT	2.58 390.805 2.63 390.935 ;
		RECT	3.84 390.805 3.89 390.935 ;
		RECT	5.675 390.805 5.725 390.935 ;
		RECT	3.06 391.035 3.11 391.165 ;
		RECT	1.085 391.495 1.135 391.625 ;
		RECT	1.405 391.535 1.455 391.585 ;
		RECT	4.47 391.535 4.6 391.585 ;
		RECT	3.06 393.455 3.11 393.585 ;
		RECT	1.57 393.685 1.62 393.815 ;
		RECT	2.58 393.685 2.63 393.815 ;
		RECT	3.84 393.685 3.89 393.815 ;
		RECT	5.675 393.685 5.725 393.815 ;
		RECT	3.06 393.915 3.11 394.045 ;
		RECT	1.085 394.375 1.135 394.505 ;
		RECT	1.405 394.415 1.455 394.465 ;
		RECT	4.47 394.415 4.6 394.465 ;
		RECT	3.06 396.335 3.11 396.465 ;
		RECT	1.57 396.565 1.62 396.695 ;
		RECT	2.58 396.565 2.63 396.695 ;
		RECT	3.84 396.565 3.89 396.695 ;
		RECT	5.675 396.565 5.725 396.695 ;
		RECT	3.06 396.795 3.11 396.925 ;
		RECT	1.085 397.255 1.135 397.385 ;
		RECT	1.405 397.295 1.455 397.345 ;
		RECT	4.47 397.295 4.6 397.345 ;
		RECT	3.06 399.215 3.11 399.345 ;
		RECT	1.57 399.445 1.62 399.575 ;
		RECT	2.58 399.445 2.63 399.575 ;
		RECT	3.84 399.445 3.89 399.575 ;
		RECT	5.675 399.445 5.725 399.575 ;
		RECT	3.06 399.675 3.11 399.805 ;
		RECT	1.085 400.135 1.135 400.265 ;
		RECT	1.405 400.175 1.455 400.225 ;
		RECT	4.47 400.175 4.6 400.225 ;
		RECT	3.06 402.095 3.11 402.225 ;
		RECT	1.57 402.325 1.62 402.455 ;
		RECT	2.58 402.325 2.63 402.455 ;
		RECT	3.84 402.325 3.89 402.455 ;
		RECT	5.675 402.325 5.725 402.455 ;
		RECT	3.06 247.035 3.11 247.165 ;
		RECT	1.085 247.495 1.135 247.625 ;
		RECT	1.405 247.535 1.455 247.585 ;
		RECT	4.47 247.535 4.6 247.585 ;
		RECT	3.06 249.455 3.11 249.585 ;
		RECT	1.57 249.685 1.62 249.815 ;
		RECT	2.58 249.685 2.63 249.815 ;
		RECT	3.84 249.685 3.89 249.815 ;
		RECT	5.675 249.685 5.725 249.815 ;
		RECT	3.06 402.555 3.11 402.685 ;
		RECT	1.085 403.015 1.135 403.145 ;
		RECT	1.405 403.055 1.455 403.105 ;
		RECT	4.47 403.055 4.6 403.105 ;
		RECT	3.06 404.975 3.11 405.105 ;
		RECT	1.57 405.205 1.62 405.335 ;
		RECT	2.58 405.205 2.63 405.335 ;
		RECT	3.84 405.205 3.89 405.335 ;
		RECT	5.675 405.205 5.725 405.335 ;
		RECT	3.06 405.435 3.11 405.565 ;
		RECT	1.085 405.895 1.135 406.025 ;
		RECT	1.405 405.935 1.455 405.985 ;
		RECT	4.47 405.935 4.6 405.985 ;
		RECT	3.06 407.855 3.11 407.985 ;
		RECT	1.57 408.085 1.62 408.215 ;
		RECT	2.58 408.085 2.63 408.215 ;
		RECT	3.84 408.085 3.89 408.215 ;
		RECT	5.675 408.085 5.725 408.215 ;
		RECT	3.06 408.315 3.11 408.445 ;
		RECT	1.085 408.775 1.135 408.905 ;
		RECT	1.405 408.815 1.455 408.865 ;
		RECT	4.47 408.815 4.6 408.865 ;
		RECT	3.06 410.735 3.11 410.865 ;
		RECT	1.57 410.965 1.62 411.095 ;
		RECT	2.58 410.965 2.63 411.095 ;
		RECT	3.84 410.965 3.89 411.095 ;
		RECT	5.675 410.965 5.725 411.095 ;
		RECT	3.06 249.915 3.11 250.045 ;
		RECT	1.085 250.375 1.135 250.505 ;
		RECT	1.405 250.415 1.455 250.465 ;
		RECT	4.47 250.415 4.6 250.465 ;
		RECT	3.06 252.335 3.11 252.465 ;
		RECT	1.57 252.565 1.62 252.695 ;
		RECT	2.58 252.565 2.63 252.695 ;
		RECT	3.84 252.565 3.89 252.695 ;
		RECT	5.675 252.565 5.725 252.695 ;
		RECT	3.06 252.795 3.11 252.925 ;
		RECT	1.085 253.255 1.135 253.385 ;
		RECT	1.405 253.295 1.455 253.345 ;
		RECT	4.47 253.295 4.6 253.345 ;
		RECT	3.06 255.215 3.11 255.345 ;
		RECT	1.57 255.445 1.62 255.575 ;
		RECT	2.58 255.445 2.63 255.575 ;
		RECT	3.84 255.445 3.89 255.575 ;
		RECT	5.675 255.445 5.725 255.575 ;
		RECT	3.06 255.675 3.11 255.805 ;
		RECT	1.085 256.135 1.135 256.265 ;
		RECT	1.405 256.175 1.455 256.225 ;
		RECT	4.47 256.175 4.6 256.225 ;
		RECT	3.06 258.095 3.11 258.225 ;
		RECT	1.57 258.325 1.62 258.455 ;
		RECT	2.58 258.325 2.63 258.455 ;
		RECT	3.84 258.325 3.89 258.455 ;
		RECT	5.675 258.325 5.725 258.455 ;
		RECT	3.06 411.195 3.11 411.325 ;
		RECT	1.085 411.655 1.135 411.785 ;
		RECT	1.405 411.695 1.455 411.745 ;
		RECT	4.47 411.695 4.6 411.745 ;
		RECT	3.06 413.615 3.11 413.745 ;
		RECT	1.57 413.845 1.62 413.975 ;
		RECT	2.58 413.845 2.63 413.975 ;
		RECT	3.84 413.845 3.89 413.975 ;
		RECT	5.675 413.845 5.725 413.975 ;
		RECT	3.06 229.755 3.11 229.885 ;
		RECT	1.085 230.215 1.135 230.345 ;
		RECT	1.405 230.255 1.455 230.305 ;
		RECT	4.47 230.255 4.6 230.305 ;
		RECT	3.06 232.175 3.11 232.305 ;
		RECT	1.57 232.405 1.62 232.535 ;
		RECT	2.58 232.405 2.63 232.535 ;
		RECT	3.84 232.405 3.89 232.535 ;
		RECT	5.675 232.405 5.725 232.535 ;
		RECT	0.435 230.215 0.485 230.345 ;
		RECT	0.435 229.755 0.485 229.885 ;
		RECT	0.435 232.175 0.485 232.305 ;
		RECT	0.435 233.095 0.485 233.225 ;
		RECT	0.435 232.635 0.485 232.765 ;
		RECT	0.435 235.055 0.485 235.185 ;
		RECT	0.435 259.015 0.485 259.145 ;
		RECT	0.435 258.555 0.485 258.685 ;
		RECT	0.435 260.975 0.485 261.105 ;
		RECT	0.435 261.895 0.485 262.025 ;
		RECT	0.435 261.435 0.485 261.565 ;
		RECT	0.435 263.855 0.485 263.985 ;
		RECT	0.435 264.775 0.485 264.905 ;
		RECT	0.435 264.315 0.485 264.445 ;
		RECT	0.435 266.735 0.485 266.865 ;
		RECT	0.435 267.655 0.485 267.785 ;
		RECT	0.435 267.195 0.485 267.325 ;
		RECT	0.435 269.615 0.485 269.745 ;
		RECT	0.435 270.535 0.485 270.665 ;
		RECT	0.435 270.075 0.485 270.205 ;
		RECT	0.435 272.495 0.485 272.625 ;
		RECT	0.435 273.415 0.485 273.545 ;
		RECT	0.435 272.955 0.485 273.085 ;
		RECT	0.435 275.375 0.485 275.505 ;
		RECT	0.435 276.295 0.485 276.425 ;
		RECT	0.435 275.835 0.485 275.965 ;
		RECT	0.435 278.255 0.485 278.385 ;
		RECT	0.435 279.175 0.485 279.305 ;
		RECT	0.435 278.715 0.485 278.845 ;
		RECT	0.435 281.135 0.485 281.265 ;
		RECT	0.435 282.055 0.485 282.185 ;
		RECT	0.435 281.595 0.485 281.725 ;
		RECT	0.435 284.015 0.485 284.145 ;
		RECT	0.435 284.935 0.485 285.065 ;
		RECT	0.435 284.475 0.485 284.605 ;
		RECT	0.435 286.895 0.485 287.025 ;
		RECT	0.435 235.975 0.485 236.105 ;
		RECT	0.435 235.515 0.485 235.645 ;
		RECT	0.435 237.935 0.485 238.065 ;
		RECT	0.435 287.815 0.485 287.945 ;
		RECT	0.435 287.355 0.485 287.485 ;
		RECT	0.435 289.775 0.485 289.905 ;
		RECT	0.435 290.695 0.485 290.825 ;
		RECT	0.435 290.235 0.485 290.365 ;
		RECT	0.435 292.655 0.485 292.785 ;
		RECT	0.435 293.575 0.485 293.705 ;
		RECT	0.435 293.115 0.485 293.245 ;
		RECT	0.435 295.535 0.485 295.665 ;
		RECT	0.435 296.455 0.485 296.585 ;
		RECT	0.435 295.995 0.485 296.125 ;
		RECT	0.435 298.415 0.485 298.545 ;
		RECT	0.435 299.335 0.485 299.465 ;
		RECT	0.435 298.875 0.485 299.005 ;
		RECT	0.435 301.295 0.485 301.425 ;
		RECT	0.435 302.215 0.485 302.345 ;
		RECT	0.435 301.755 0.485 301.885 ;
		RECT	0.435 304.175 0.485 304.305 ;
		RECT	0.435 305.095 0.485 305.225 ;
		RECT	0.435 304.635 0.485 304.765 ;
		RECT	0.435 307.055 0.485 307.185 ;
		RECT	0.435 307.975 0.485 308.105 ;
		RECT	0.435 307.515 0.485 307.645 ;
		RECT	0.435 309.935 0.485 310.065 ;
		RECT	0.435 310.855 0.485 310.985 ;
		RECT	0.435 310.395 0.485 310.525 ;
		RECT	0.435 312.815 0.485 312.945 ;
		RECT	0.435 313.735 0.485 313.865 ;
		RECT	0.435 313.275 0.485 313.405 ;
		RECT	0.435 315.695 0.485 315.825 ;
		RECT	0.435 238.855 0.485 238.985 ;
		RECT	0.435 238.395 0.485 238.525 ;
		RECT	0.435 240.815 0.485 240.945 ;
		RECT	0.435 316.615 0.485 316.745 ;
		RECT	0.435 316.155 0.485 316.285 ;
		RECT	0.435 318.575 0.485 318.705 ;
		RECT	0.435 319.495 0.485 319.625 ;
		RECT	0.435 319.035 0.485 319.165 ;
		RECT	0.435 321.455 0.485 321.585 ;
		RECT	0.435 322.375 0.485 322.505 ;
		RECT	0.435 321.915 0.485 322.045 ;
		RECT	0.435 324.335 0.485 324.465 ;
		RECT	0.435 325.255 0.485 325.385 ;
		RECT	0.435 324.795 0.485 324.925 ;
		RECT	0.435 327.215 0.485 327.345 ;
		RECT	0.435 328.135 0.485 328.265 ;
		RECT	0.435 327.675 0.485 327.805 ;
		RECT	0.435 330.095 0.485 330.225 ;
		RECT	0.435 331.015 0.485 331.145 ;
		RECT	0.435 330.555 0.485 330.685 ;
		RECT	0.435 332.975 0.485 333.105 ;
		RECT	0.435 333.895 0.485 334.025 ;
		RECT	0.435 333.435 0.485 333.565 ;
		RECT	0.435 335.855 0.485 335.985 ;
		RECT	0.435 336.775 0.485 336.905 ;
		RECT	0.435 336.315 0.485 336.445 ;
		RECT	0.435 338.735 0.485 338.865 ;
		RECT	0.435 339.655 0.485 339.785 ;
		RECT	0.435 339.195 0.485 339.325 ;
		RECT	0.435 341.615 0.485 341.745 ;
		RECT	0.435 342.535 0.485 342.665 ;
		RECT	0.435 342.075 0.485 342.205 ;
		RECT	0.435 344.495 0.485 344.625 ;
		RECT	0.435 241.735 0.485 241.865 ;
		RECT	0.435 241.275 0.485 241.405 ;
		RECT	0.435 243.695 0.485 243.825 ;
		RECT	0.435 345.415 0.485 345.545 ;
		RECT	0.435 344.955 0.485 345.085 ;
		RECT	0.435 347.375 0.485 347.505 ;
		RECT	0.435 348.295 0.485 348.425 ;
		RECT	0.435 347.835 0.485 347.965 ;
		RECT	0.435 350.255 0.485 350.385 ;
		RECT	0.435 351.175 0.485 351.305 ;
		RECT	0.435 350.715 0.485 350.845 ;
		RECT	0.435 353.135 0.485 353.265 ;
		RECT	0.435 354.055 0.485 354.185 ;
		RECT	0.435 353.595 0.485 353.725 ;
		RECT	0.435 356.015 0.485 356.145 ;
		RECT	0.435 356.935 0.485 357.065 ;
		RECT	0.435 356.475 0.485 356.605 ;
		RECT	0.435 358.895 0.485 359.025 ;
		RECT	0.435 359.815 0.485 359.945 ;
		RECT	0.435 359.355 0.485 359.485 ;
		RECT	0.435 361.775 0.485 361.905 ;
		RECT	0.435 362.695 0.485 362.825 ;
		RECT	0.435 362.235 0.485 362.365 ;
		RECT	0.435 364.655 0.485 364.785 ;
		RECT	0.435 365.575 0.485 365.705 ;
		RECT	0.435 365.115 0.485 365.245 ;
		RECT	0.435 367.535 0.485 367.665 ;
		RECT	0.435 368.455 0.485 368.585 ;
		RECT	0.435 367.995 0.485 368.125 ;
		RECT	0.435 370.415 0.485 370.545 ;
		RECT	0.435 371.335 0.485 371.465 ;
		RECT	0.435 370.875 0.485 371.005 ;
		RECT	0.435 373.295 0.485 373.425 ;
		RECT	0.435 244.615 0.485 244.745 ;
		RECT	0.435 244.155 0.485 244.285 ;
		RECT	0.435 246.575 0.485 246.705 ;
		RECT	0.435 374.215 0.485 374.345 ;
		RECT	0.435 373.755 0.485 373.885 ;
		RECT	0.435 376.175 0.485 376.305 ;
		RECT	0.435 377.095 0.485 377.225 ;
		RECT	0.435 376.635 0.485 376.765 ;
		RECT	0.435 379.055 0.485 379.185 ;
		RECT	0.435 379.975 0.485 380.105 ;
		RECT	0.435 379.515 0.485 379.645 ;
		RECT	0.435 381.935 0.485 382.065 ;
		RECT	0.435 382.855 0.485 382.985 ;
		RECT	0.435 382.395 0.485 382.525 ;
		RECT	0.435 384.815 0.485 384.945 ;
		RECT	0.435 385.735 0.485 385.865 ;
		RECT	0.435 385.275 0.485 385.405 ;
		RECT	0.435 387.695 0.485 387.825 ;
		RECT	0.435 388.615 0.485 388.745 ;
		RECT	0.435 388.155 0.485 388.285 ;
		RECT	0.435 390.575 0.485 390.705 ;
		RECT	0.435 391.495 0.485 391.625 ;
		RECT	0.435 391.035 0.485 391.165 ;
		RECT	0.435 393.455 0.485 393.585 ;
		RECT	0.435 394.375 0.485 394.505 ;
		RECT	0.435 393.915 0.485 394.045 ;
		RECT	0.435 396.335 0.485 396.465 ;
		RECT	0.435 397.255 0.485 397.385 ;
		RECT	0.435 396.795 0.485 396.925 ;
		RECT	0.435 399.215 0.485 399.345 ;
		RECT	0.435 400.135 0.485 400.265 ;
		RECT	0.435 399.675 0.485 399.805 ;
		RECT	0.435 402.095 0.485 402.225 ;
		RECT	0.435 247.495 0.485 247.625 ;
		RECT	0.435 247.035 0.485 247.165 ;
		RECT	0.435 249.455 0.485 249.585 ;
		RECT	0.435 403.015 0.485 403.145 ;
		RECT	0.435 402.555 0.485 402.685 ;
		RECT	0.435 404.975 0.485 405.105 ;
		RECT	0.435 405.895 0.485 406.025 ;
		RECT	0.435 405.435 0.485 405.565 ;
		RECT	0.435 407.855 0.485 407.985 ;
		RECT	0.435 408.775 0.485 408.905 ;
		RECT	0.435 408.315 0.485 408.445 ;
		RECT	0.435 410.735 0.485 410.865 ;
		RECT	0.435 411.655 0.485 411.785 ;
		RECT	0.435 411.195 0.485 411.325 ;
		RECT	0.435 413.615 0.485 413.745 ;
		RECT	0.435 250.375 0.485 250.505 ;
		RECT	0.435 249.915 0.485 250.045 ;
		RECT	0.435 252.335 0.485 252.465 ;
		RECT	0.435 253.255 0.485 253.385 ;
		RECT	0.435 252.795 0.485 252.925 ;
		RECT	0.435 255.215 0.485 255.345 ;
		RECT	0.435 256.135 0.485 256.265 ;
		RECT	0.435 255.675 0.485 255.805 ;
		RECT	0.435 258.095 0.485 258.225 ;
		RECT	20.085 186.875 20.265 187.005 ;
		RECT	20.08 192.86 20.21 193.04 ;
		RECT	20.08 221.89 20.21 222.07 ;
		RECT	20.085 227.855 20.265 227.985 ;
		RECT	20.395 188.455 20.575 188.585 ;
		RECT	20.53 190.46 20.58 190.59 ;
		RECT	20.53 193.375 20.58 193.505 ;
		RECT	20.53 194.36 20.58 194.49 ;
		RECT	20.53 196.33 20.58 196.46 ;
		RECT	20.53 197.31 20.58 197.44 ;
		RECT	20.53 198.295 20.58 198.425 ;
		RECT	20.53 201.25 20.58 201.38 ;
		RECT	20.53 208.63 20.58 208.76 ;
		RECT	20.53 209.61 20.58 209.74 ;
		RECT	20.53 213.55 20.58 213.68 ;
		RECT	20.53 216.5 20.58 216.63 ;
		RECT	20.53 217.485 20.58 217.615 ;
		RECT	20.53 218.47 20.58 218.6 ;
		RECT	20.53 220.435 20.58 220.565 ;
		RECT	20.53 221.42 20.58 221.55 ;
		RECT	20.53 224.34 20.58 224.47 ;
		RECT	20.395 226.34 20.575 226.47 ;
		RECT	20.875 187.105 21.055 187.235 ;
		RECT	20.875 227.625 21.055 227.755 ;
		RECT	20.085 187.58 20.265 187.71 ;
		RECT	20.11 227.12 20.24 227.3 ;
		RECT	20.12 189.915 20.17 190.045 ;
		RECT	20.12 193.87 20.17 194 ;
		RECT	20.12 197.805 20.17 197.935 ;
		RECT	20.12 201.74 20.17 201.87 ;
		RECT	20.12 205.675 20.17 205.805 ;
		RECT	20.12 209.12 20.17 209.25 ;
		RECT	20.12 213.055 20.17 213.185 ;
		RECT	20.12 216.995 20.17 217.125 ;
		RECT	20.12 220.93 20.17 221.06 ;
		RECT	20.12 224.88 20.17 225.01 ;
		RECT	14.965 186.875 15.015 187.005 ;
		RECT	19.485 186.875 19.535 187.005 ;
		RECT	14.765 186.875 14.815 187.005 ;
		RECT	19.685 186.875 19.735 187.005 ;
		RECT	14.965 227.855 15.015 227.985 ;
		RECT	19.485 227.855 19.535 227.985 ;
		RECT	14.765 227.855 14.815 227.985 ;
		RECT	19.685 227.855 19.735 227.985 ;
		RECT	20.395 186.645 20.575 186.775 ;
		RECT	20.7 187.105 20.75 187.235 ;
		RECT	20.085 187.965 20.265 188.095 ;
		RECT	20.9 188.74 21.03 188.79 ;
		RECT	20.085 188.945 20.265 189.075 ;
		RECT	20.39 189.44 20.44 189.57 ;
		RECT	20.9 189.72 21.03 189.77 ;
		RECT	20.685 190.19 20.735 190.32 ;
		RECT	20.335 190.19 20.385 190.32 ;
		RECT	20.12 190.915 20.17 191.045 ;
		RECT	20.875 191.41 21.055 191.54 ;
		RECT	20.12 191.9 20.17 192.03 ;
		RECT	20.08 192.185 20.21 192.235 ;
		RECT	20.875 192.39 21.055 192.52 ;
		RECT	20.12 194.855 20.17 194.985 ;
		RECT	20.875 195.345 21.055 195.475 ;
		RECT	20.12 195.835 20.17 195.965 ;
		RECT	20.12 196.82 20.17 196.95 ;
		RECT	20.12 198.79 20.17 198.92 ;
		RECT	20.875 199.28 21.055 199.41 ;
		RECT	20.12 199.77 20.17 199.9 ;
		RECT	20.875 200.265 21.055 200.395 ;
		RECT	20.12 200.755 20.17 200.885 ;
		RECT	20.53 202.235 20.58 202.365 ;
		RECT	20.12 202.73 20.17 202.86 ;
		RECT	20.875 203.215 21.055 203.345 ;
		RECT	20.12 203.71 20.17 203.84 ;
		RECT	20.505 204.185 20.555 204.315 ;
		RECT	20.685 204.495 20.735 204.625 ;
		RECT	20.335 204.495 20.385 204.625 ;
		RECT	20.345 204.81 20.395 204.94 ;
		RECT	20.9 205.47 21.03 205.52 ;
		RECT	20.9 205.965 21.03 206.015 ;
		RECT	20.12 206.66 20.17 206.79 ;
		RECT	20.875 207.15 21.055 207.28 ;
		RECT	20.875 207.645 21.055 207.775 ;
		RECT	20.12 208.135 20.17 208.265 ;
		RECT	20.9 208.915 21.03 208.965 ;
		RECT	20.9 209.405 21.03 209.455 ;
		RECT	20.345 209.925 20.395 210.055 ;
		RECT	20.685 210.27 20.735 210.4 ;
		RECT	20.335 210.27 20.385 210.4 ;
		RECT	20.12 211.085 20.17 211.215 ;
		RECT	20.875 211.58 21.055 211.71 ;
		RECT	20.12 212.075 20.17 212.205 ;
		RECT	20.53 212.565 20.58 212.695 ;
		RECT	20.12 214.04 20.17 214.17 ;
		RECT	20.875 214.535 21.055 214.665 ;
		RECT	20.12 215.025 20.17 215.155 ;
		RECT	20.875 215.515 21.055 215.645 ;
		RECT	20.12 216.01 20.17 216.14 ;
		RECT	20.12 217.975 20.17 218.105 ;
		RECT	20.12 218.96 20.17 219.09 ;
		RECT	20.875 219.455 21.055 219.585 ;
		RECT	20.12 219.945 20.17 220.075 ;
		RECT	20.08 220.72 20.21 220.77 ;
		RECT	20.08 222.2 20.21 222.25 ;
		RECT	20.875 222.405 21.055 222.535 ;
		RECT	20.08 222.69 20.21 222.74 ;
		RECT	20.12 222.895 20.17 223.025 ;
		RECT	20.875 223.355 21.055 223.485 ;
		RECT	20.12 223.88 20.17 224.01 ;
		RECT	20.685 224.61 20.735 224.74 ;
		RECT	20.335 224.61 20.385 224.74 ;
		RECT	20.9 225.155 21.03 225.205 ;
		RECT	20.39 225.355 20.44 225.485 ;
		RECT	20.085 225.85 20.265 225.98 ;
		RECT	20.9 226.135 21.03 226.185 ;
		RECT	20.085 226.835 20.265 226.965 ;
		RECT	20.7 227.625 20.75 227.755 ;
		RECT	20.395 228.085 20.575 228.215 ;
		RECT	14.965 187.58 15.015 187.71 ;
		RECT	14.99 190.915 15.04 191.045 ;
		RECT	14.99 191.9 15.04 192.03 ;
		RECT	14.99 192.185 15.04 192.235 ;
		RECT	14.99 194.855 15.04 194.985 ;
		RECT	14.99 195.835 15.04 195.965 ;
		RECT	14.99 196.82 15.04 196.95 ;
		RECT	14.99 198.79 15.04 198.92 ;
		RECT	14.99 199.77 15.04 199.9 ;
		RECT	14.99 200.755 15.04 200.885 ;
		RECT	14.99 202.73 15.04 202.86 ;
		RECT	14.99 203.71 15.04 203.84 ;
		RECT	14.965 206.66 15.015 206.79 ;
		RECT	14.965 208.135 15.015 208.265 ;
		RECT	14.99 211.085 15.04 211.215 ;
		RECT	14.99 212.075 15.04 212.205 ;
		RECT	14.99 214.04 15.04 214.17 ;
		RECT	14.99 215.025 15.04 215.155 ;
		RECT	14.99 216.01 15.04 216.14 ;
		RECT	14.99 217.975 15.04 218.105 ;
		RECT	14.99 218.96 15.04 219.09 ;
		RECT	14.99 219.945 15.04 220.075 ;
		RECT	14.99 220.72 15.04 220.77 ;
		RECT	14.99 222.895 15.04 223.025 ;
		RECT	14.99 223.88 15.04 224.01 ;
		RECT	14.965 227.145 15.015 227.275 ;
		RECT	19.485 187.58 19.535 187.71 ;
		RECT	19.465 201.715 19.595 201.895 ;
		RECT	19.465 213.03 19.595 213.21 ;
		RECT	19.465 220.905 19.595 221.085 ;
		RECT	19.485 227.145 19.535 227.275 ;
		RECT	19.875 204.185 19.925 204.315 ;
		RECT	19.875 210.61 19.925 210.74 ;
		RECT	19.7 187.965 19.75 188.095 ;
		RECT	19.7 188.945 19.75 189.075 ;
		RECT	19.7 190.915 19.75 191.045 ;
		RECT	19.7 191.9 19.75 192.03 ;
		RECT	19.7 192.185 19.75 192.235 ;
		RECT	19.7 194.855 19.75 194.985 ;
		RECT	19.7 195.835 19.75 195.965 ;
		RECT	19.7 196.82 19.75 196.95 ;
		RECT	19.7 198.79 19.75 198.92 ;
		RECT	19.7 199.77 19.75 199.9 ;
		RECT	19.7 200.755 19.75 200.885 ;
		RECT	19.7 202.73 19.75 202.86 ;
		RECT	19.7 203.71 19.75 203.84 ;
		RECT	19.7 206.66 19.75 206.79 ;
		RECT	19.7 208.135 19.75 208.265 ;
		RECT	19.7 211.085 19.75 211.215 ;
		RECT	19.7 212.075 19.75 212.205 ;
		RECT	19.7 214.04 19.75 214.17 ;
		RECT	19.7 215.025 19.75 215.155 ;
		RECT	19.7 216.01 19.75 216.14 ;
		RECT	19.7 217.975 19.75 218.105 ;
		RECT	19.7 218.96 19.75 219.09 ;
		RECT	19.7 219.945 19.75 220.075 ;
		RECT	19.7 220.72 19.75 220.77 ;
		RECT	19.465 221.89 19.595 222.07 ;
		RECT	19.7 222.895 19.75 223.025 ;
		RECT	19.7 223.88 19.75 224.01 ;
		RECT	19.7 225.85 19.75 225.98 ;
		RECT	19.7 226.835 19.75 226.965 ;
		RECT	14.765 187.965 14.815 188.095 ;
		RECT	14.765 188.945 14.815 189.075 ;
		RECT	14.74 190.915 14.79 191.045 ;
		RECT	14.74 191.9 14.79 192.03 ;
		RECT	14.74 192.185 14.79 192.235 ;
		RECT	14.74 194.855 14.79 194.985 ;
		RECT	14.74 195.835 14.79 195.965 ;
		RECT	14.74 196.82 14.79 196.95 ;
		RECT	14.74 198.79 14.79 198.92 ;
		RECT	14.74 199.77 14.79 199.9 ;
		RECT	14.74 200.755 14.79 200.885 ;
		RECT	14.74 202.73 14.79 202.86 ;
		RECT	14.74 203.71 14.79 203.84 ;
		RECT	14.765 206.66 14.815 206.79 ;
		RECT	14.765 208.135 14.815 208.265 ;
		RECT	14.74 211.085 14.79 211.215 ;
		RECT	14.74 212.075 14.79 212.205 ;
		RECT	14.74 214.04 14.79 214.17 ;
		RECT	14.74 215.025 14.79 215.155 ;
		RECT	14.74 216.01 14.79 216.14 ;
		RECT	14.74 217.975 14.79 218.105 ;
		RECT	14.74 218.96 14.79 219.09 ;
		RECT	14.74 219.945 14.79 220.075 ;
		RECT	14.74 220.72 14.79 220.77 ;
		RECT	14.74 222.895 14.79 223.025 ;
		RECT	14.74 223.88 14.79 224.01 ;
		RECT	14.765 225.85 14.815 225.98 ;
		RECT	14.765 226.835 14.815 226.965 ;
		RECT	14.565 204.185 14.615 204.315 ;
		RECT	14.565 210.61 14.615 210.74 ;
		RECT	14.965 187.965 15.015 188.095 ;
		RECT	15.335 187.965 15.385 188.095 ;
		RECT	15.875 187.965 15.925 188.095 ;
		RECT	16.415 187.965 16.465 188.095 ;
		RECT	16.955 187.965 17.005 188.095 ;
		RECT	17.495 187.965 17.545 188.095 ;
		RECT	18.035 187.965 18.085 188.095 ;
		RECT	18.575 187.965 18.625 188.095 ;
		RECT	19.115 187.965 19.165 188.095 ;
		RECT	14.565 188.74 14.615 188.79 ;
		RECT	14.965 188.945 15.015 189.075 ;
		RECT	15.335 189.44 15.385 189.57 ;
		RECT	15.875 189.44 15.925 189.57 ;
		RECT	16.415 189.44 16.465 189.57 ;
		RECT	16.955 189.44 17.005 189.57 ;
		RECT	17.495 189.44 17.545 189.57 ;
		RECT	18.035 189.44 18.085 189.57 ;
		RECT	18.575 189.44 18.625 189.57 ;
		RECT	19.115 189.44 19.165 189.57 ;
		RECT	14.565 189.72 14.615 189.77 ;
		RECT	14.99 189.915 15.04 190.045 ;
		RECT	14.865 190.19 14.915 190.32 ;
		RECT	15.335 190.19 15.385 190.32 ;
		RECT	15.875 190.19 15.925 190.32 ;
		RECT	16.415 190.19 16.465 190.32 ;
		RECT	16.955 190.19 17.005 190.32 ;
		RECT	17.495 190.19 17.545 190.32 ;
		RECT	18.035 190.19 18.085 190.32 ;
		RECT	18.575 190.19 18.625 190.32 ;
		RECT	19.115 190.19 19.165 190.32 ;
		RECT	14.565 191.41 14.615 191.54 ;
		RECT	14.565 192.39 14.615 192.52 ;
		RECT	14.745 192.885 14.795 193.015 ;
		RECT	14.99 193.87 15.04 194 ;
		RECT	14.565 195.345 14.615 195.475 ;
		RECT	14.99 197.805 15.04 197.935 ;
		RECT	14.565 199.255 14.615 199.435 ;
		RECT	14.565 200.24 14.615 200.425 ;
		RECT	14.99 201.715 15.04 201.895 ;
		RECT	14.565 203.19 14.615 203.37 ;
		RECT	13.8 204.185 13.85 204.315 ;
		RECT	14.865 204.495 14.915 204.625 ;
		RECT	15.335 204.495 15.385 204.625 ;
		RECT	15.875 204.495 15.925 204.625 ;
		RECT	16.415 204.495 16.465 204.625 ;
		RECT	16.955 204.495 17.005 204.625 ;
		RECT	17.495 204.495 17.545 204.625 ;
		RECT	18.035 204.495 18.085 204.625 ;
		RECT	18.575 204.495 18.625 204.625 ;
		RECT	19.115 204.495 19.165 204.625 ;
		RECT	15.335 204.81 15.385 204.94 ;
		RECT	15.875 204.81 15.925 204.94 ;
		RECT	16.415 204.81 16.465 204.94 ;
		RECT	16.955 204.81 17.005 204.94 ;
		RECT	17.495 204.81 17.545 204.94 ;
		RECT	18.035 204.81 18.085 204.94 ;
		RECT	18.575 204.81 18.625 204.94 ;
		RECT	19.115 204.81 19.165 204.94 ;
		RECT	14.565 205.47 14.615 205.52 ;
		RECT	14.965 205.675 15.015 205.805 ;
		RECT	14.565 205.965 14.615 206.015 ;
		RECT	15.335 206.66 15.385 206.79 ;
		RECT	15.875 206.66 15.925 206.79 ;
		RECT	16.415 206.66 16.465 206.79 ;
		RECT	16.955 206.66 17.005 206.79 ;
		RECT	17.495 206.66 17.545 206.79 ;
		RECT	18.035 206.66 18.085 206.79 ;
		RECT	18.575 206.66 18.625 206.79 ;
		RECT	19.115 206.66 19.165 206.79 ;
		RECT	14.565 207.12 14.615 207.31 ;
		RECT	14.565 207.615 14.615 207.805 ;
		RECT	15.335 208.135 15.385 208.265 ;
		RECT	15.875 208.135 15.925 208.265 ;
		RECT	16.415 208.135 16.465 208.265 ;
		RECT	16.955 208.135 17.005 208.265 ;
		RECT	17.495 208.135 17.545 208.265 ;
		RECT	18.035 208.135 18.085 208.265 ;
		RECT	18.575 208.135 18.625 208.265 ;
		RECT	19.115 208.135 19.165 208.265 ;
		RECT	14.565 208.915 14.615 208.965 ;
		RECT	14.965 209.12 15.015 209.25 ;
		RECT	14.565 209.405 14.615 209.455 ;
		RECT	15.335 209.925 15.385 210.055 ;
		RECT	15.875 209.925 15.925 210.055 ;
		RECT	16.415 209.925 16.465 210.055 ;
		RECT	16.955 209.925 17.005 210.055 ;
		RECT	17.495 209.925 17.545 210.055 ;
		RECT	18.035 209.925 18.085 210.055 ;
		RECT	18.575 209.925 18.625 210.055 ;
		RECT	19.115 209.925 19.165 210.055 ;
		RECT	14.865 210.27 14.915 210.4 ;
		RECT	15.335 210.27 15.385 210.4 ;
		RECT	15.875 210.27 15.925 210.4 ;
		RECT	16.415 210.27 16.465 210.4 ;
		RECT	16.955 210.27 17.005 210.4 ;
		RECT	17.495 210.27 17.545 210.4 ;
		RECT	18.035 210.27 18.085 210.4 ;
		RECT	18.575 210.27 18.625 210.4 ;
		RECT	19.115 210.27 19.165 210.4 ;
		RECT	13.8 210.61 13.85 210.74 ;
		RECT	14.565 211.555 14.615 211.735 ;
		RECT	14.99 213.03 15.04 213.21 ;
		RECT	14.565 214.505 14.615 214.69 ;
		RECT	14.565 215.49 14.615 215.67 ;
		RECT	14.99 216.97 15.04 217.15 ;
		RECT	14.565 219.43 14.615 219.61 ;
		RECT	14.99 220.93 15.04 221.06 ;
		RECT	14.745 221.915 14.795 222.045 ;
		RECT	14.565 222.405 14.615 222.535 ;
		RECT	14.565 223.33 14.615 223.51 ;
		RECT	14.865 224.61 14.915 224.74 ;
		RECT	15.335 224.61 15.385 224.74 ;
		RECT	15.875 224.61 15.925 224.74 ;
		RECT	16.415 224.61 16.465 224.74 ;
		RECT	16.955 224.61 17.005 224.74 ;
		RECT	17.495 224.61 17.545 224.74 ;
		RECT	18.035 224.61 18.085 224.74 ;
		RECT	18.575 224.61 18.625 224.74 ;
		RECT	19.115 224.61 19.165 224.74 ;
		RECT	14.99 224.88 15.04 225.01 ;
		RECT	14.565 225.155 14.615 225.205 ;
		RECT	15.335 225.355 15.385 225.485 ;
		RECT	15.875 225.355 15.925 225.485 ;
		RECT	16.415 225.355 16.465 225.485 ;
		RECT	16.955 225.355 17.005 225.485 ;
		RECT	17.495 225.355 17.545 225.485 ;
		RECT	18.035 225.355 18.085 225.485 ;
		RECT	18.575 225.355 18.625 225.485 ;
		RECT	19.115 225.355 19.165 225.485 ;
		RECT	14.965 225.85 15.015 225.98 ;
		RECT	14.565 226.135 14.615 226.185 ;
		RECT	14.965 226.835 15.015 226.965 ;
		RECT	15.335 226.835 15.385 226.965 ;
		RECT	15.875 226.835 15.925 226.965 ;
		RECT	16.415 226.835 16.465 226.965 ;
		RECT	16.955 226.835 17.005 226.965 ;
		RECT	17.495 226.835 17.545 226.965 ;
		RECT	18.035 226.835 18.085 226.965 ;
		RECT	18.575 226.835 18.625 226.965 ;
		RECT	19.115 226.835 19.165 226.965 ;
		RECT	19.465 187.94 19.595 188.12 ;
		RECT	19.85 188.74 19.98 188.79 ;
		RECT	19.465 188.985 19.595 189.035 ;
		RECT	19.85 189.72 19.98 189.77 ;
		RECT	19.465 190.89 19.595 191.07 ;
		RECT	19.885 191.41 19.935 191.54 ;
		RECT	19.465 191.94 19.595 191.99 ;
		RECT	19.465 192.185 19.595 192.235 ;
		RECT	19.885 192.39 19.935 192.52 ;
		RECT	19.7 192.885 19.75 193.015 ;
		RECT	19.465 194.83 19.595 195.01 ;
		RECT	19.885 195.345 19.935 195.475 ;
		RECT	19.465 195.81 19.595 195.99 ;
		RECT	19.465 196.795 19.595 196.975 ;
		RECT	19.465 198.765 19.595 198.945 ;
		RECT	19.885 199.28 19.935 199.41 ;
		RECT	19.465 199.745 19.595 199.925 ;
		RECT	19.885 200.265 19.935 200.395 ;
		RECT	19.465 200.73 19.595 200.91 ;
		RECT	19.465 202.705 19.595 202.885 ;
		RECT	19.885 203.215 19.935 203.345 ;
		RECT	19.465 203.685 19.595 203.865 ;
		RECT	19.85 205.47 19.98 205.52 ;
		RECT	19.85 205.965 19.98 206.015 ;
		RECT	19.465 206.635 19.595 206.815 ;
		RECT	19.885 207.15 19.935 207.28 ;
		RECT	19.885 207.645 19.935 207.775 ;
		RECT	19.465 208.11 19.595 208.29 ;
		RECT	19.85 208.915 19.98 208.965 ;
		RECT	19.85 209.405 19.98 209.455 ;
		RECT	19.465 211.06 19.595 211.24 ;
		RECT	19.885 211.58 19.935 211.71 ;
		RECT	19.465 212.05 19.595 212.23 ;
		RECT	19.465 214.015 19.595 214.195 ;
		RECT	19.885 214.535 19.935 214.665 ;
		RECT	19.465 215 19.595 215.18 ;
		RECT	19.885 215.515 19.935 215.645 ;
		RECT	19.465 215.985 19.595 216.165 ;
		RECT	19.465 217.95 19.595 218.13 ;
		RECT	19.465 218.935 19.595 219.115 ;
		RECT	19.885 219.455 19.935 219.585 ;
		RECT	19.465 219.92 19.595 220.1 ;
		RECT	19.465 220.72 19.595 220.77 ;
		RECT	19.7 221.915 19.75 222.045 ;
		RECT	19.885 222.405 19.935 222.535 ;
		RECT	19.465 222.87 19.595 223.05 ;
		RECT	19.885 223.355 19.935 223.485 ;
		RECT	19.465 223.855 19.595 224.035 ;
		RECT	19.85 225.155 19.98 225.205 ;
		RECT	19.465 225.89 19.595 225.94 ;
		RECT	19.885 226.135 19.935 226.185 ;
		RECT	19.465 226.875 19.595 226.925 ;
	END

END rf2_32x128_wm1

END LIBRARY

